magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< error_p >>
rect 22800 4869 22806 4875
rect 22797 4863 22800 4869
<< metal1 >>
rect 0 44952 200 45152
rect 28872 44952 29072 45152
rect 7722 41626 7780 41632
rect 7780 41568 7892 41626
rect 8050 41623 8102 41629
rect 7722 41562 7780 41568
rect 8050 41565 8102 41571
rect 8350 41623 8402 41629
rect 8350 41565 8402 41571
rect 8650 41623 8702 41629
rect 8650 41565 8702 41571
rect 8950 41623 9002 41629
rect 8950 41565 9002 41571
rect 9250 41623 9302 41629
rect 9250 41565 9302 41571
rect 9550 41623 9602 41629
rect 9550 41565 9602 41571
rect 9850 41623 9902 41629
rect 9850 41565 9902 41571
rect 10150 41626 10202 41629
rect 10278 41626 10336 41632
rect 10150 41623 10278 41626
rect 10202 41571 10278 41623
rect 10150 41568 10278 41571
rect 10150 41565 10202 41568
rect 10278 41562 10336 41568
rect 12922 41626 12980 41632
rect 12980 41568 13092 41626
rect 13250 41623 13302 41629
rect 12922 41562 12980 41568
rect 13250 41565 13302 41571
rect 13550 41623 13602 41629
rect 13550 41565 13602 41571
rect 13850 41623 13902 41629
rect 13850 41565 13902 41571
rect 14150 41623 14202 41629
rect 14150 41565 14202 41571
rect 14450 41623 14502 41629
rect 14450 41565 14502 41571
rect 14750 41623 14802 41629
rect 14750 41565 14802 41571
rect 15050 41623 15102 41629
rect 15050 41565 15102 41571
rect 15350 41626 15402 41629
rect 15478 41626 15536 41632
rect 15350 41623 15478 41626
rect 15402 41571 15478 41623
rect 15350 41568 15478 41571
rect 15350 41565 15402 41568
rect 15478 41562 15536 41568
rect 2664 41342 2724 41348
rect 2664 41276 2724 41282
rect 2964 41342 3024 41348
rect 2964 41276 3024 41282
rect 3264 41342 3324 41348
rect 3264 41276 3324 41282
rect 3564 41342 3624 41348
rect 3564 41276 3624 41282
rect 3864 41342 3924 41348
rect 3864 41276 3924 41282
rect 4164 41342 4224 41348
rect 4164 41276 4224 41282
rect 4464 41342 4524 41348
rect 4464 41276 4524 41282
rect 4764 41342 4824 41348
rect 4764 41276 4824 41282
rect 21352 41325 21410 41331
rect 21453 41325 21505 41328
rect 21410 41322 21505 41325
rect 21410 41270 21453 41322
rect 21410 41267 21505 41270
rect 21352 41261 21410 41267
rect 21453 41264 21505 41267
rect 21753 41322 21805 41328
rect 21753 41264 21805 41270
rect 22053 41322 22105 41328
rect 22053 41264 22105 41270
rect 22353 41322 22405 41328
rect 22353 41264 22405 41270
rect 22653 41322 22705 41328
rect 22653 41264 22705 41270
rect 22953 41322 23005 41328
rect 22953 41264 23005 41270
rect 23253 41322 23305 41328
rect 23253 41264 23305 41270
rect 23553 41322 23605 41328
rect 23858 41325 23916 41331
rect 23553 41264 23605 41270
rect 23776 41267 23858 41325
rect 23858 41261 23916 41267
rect 7745 40500 7815 40506
rect 10252 40500 10322 40506
rect 7815 40436 7892 40494
rect 10176 40436 10252 40494
rect 7745 40424 7815 40430
rect 10252 40424 10322 40430
rect 12945 40500 13015 40506
rect 15452 40500 15522 40506
rect 13015 40436 13092 40494
rect 15376 40436 15452 40494
rect 12945 40424 13015 40430
rect 15452 40424 15522 40430
rect 7716 40290 7786 40296
rect 10272 40290 10342 40296
rect 7786 40226 7892 40284
rect 10176 40226 10272 40284
rect 7716 40214 7786 40220
rect 10272 40214 10342 40220
rect 12916 40290 12986 40296
rect 15472 40290 15542 40296
rect 12986 40226 13092 40284
rect 15376 40226 15472 40284
rect 12916 40214 12986 40220
rect 15472 40214 15542 40220
rect 2667 40206 2719 40212
rect 2667 40148 2719 40154
rect 2967 40206 3019 40212
rect 2967 40148 3019 40154
rect 3267 40206 3319 40212
rect 3267 40148 3319 40154
rect 3567 40206 3619 40212
rect 3567 40148 3619 40154
rect 3867 40206 3919 40212
rect 3867 40148 3919 40154
rect 4167 40206 4219 40212
rect 4167 40148 4219 40154
rect 4467 40206 4519 40212
rect 4467 40148 4519 40154
rect 4767 40206 4819 40212
rect 21467 40193 21519 40196
rect 4767 40148 4819 40154
rect 21326 40135 21332 40193
rect 21390 40190 21519 40193
rect 21390 40138 21467 40190
rect 21390 40135 21519 40138
rect 21467 40132 21519 40135
rect 21767 40190 21819 40196
rect 21767 40132 21819 40138
rect 22067 40190 22119 40196
rect 22067 40132 22119 40138
rect 22367 40190 22419 40196
rect 22367 40132 22419 40138
rect 22667 40190 22719 40196
rect 22667 40132 22719 40138
rect 22967 40190 23019 40196
rect 22967 40132 23019 40138
rect 23267 40190 23319 40196
rect 23267 40132 23319 40138
rect 23567 40190 23619 40196
rect 23888 40193 23946 40199
rect 23567 40132 23619 40138
rect 23776 40135 23888 40193
rect 23888 40129 23946 40135
rect 7752 39152 7810 39158
rect 7810 39094 7892 39152
rect 8049 39149 8101 39155
rect 7752 39088 7810 39094
rect 8049 39091 8101 39097
rect 8349 39149 8401 39155
rect 8349 39091 8401 39097
rect 8649 39149 8701 39155
rect 8649 39091 8701 39097
rect 8949 39149 9001 39155
rect 8949 39091 9001 39097
rect 9249 39149 9301 39155
rect 9249 39091 9301 39097
rect 9549 39149 9601 39155
rect 9549 39091 9601 39097
rect 9849 39149 9901 39155
rect 9849 39091 9901 39097
rect 10149 39152 10201 39155
rect 10258 39152 10316 39158
rect 10149 39149 10258 39152
rect 10201 39097 10258 39149
rect 10149 39094 10258 39097
rect 10149 39091 10201 39094
rect 10258 39088 10316 39094
rect 12952 39152 13010 39158
rect 13010 39094 13092 39152
rect 13249 39149 13301 39155
rect 12952 39088 13010 39094
rect 13249 39091 13301 39097
rect 13549 39149 13601 39155
rect 13549 39091 13601 39097
rect 13849 39149 13901 39155
rect 13849 39091 13901 39097
rect 14149 39149 14201 39155
rect 14149 39091 14201 39097
rect 14449 39149 14501 39155
rect 14449 39091 14501 39097
rect 14749 39149 14801 39155
rect 14749 39091 14801 39097
rect 15049 39149 15101 39155
rect 15049 39091 15101 39097
rect 15349 39152 15401 39155
rect 15458 39152 15516 39158
rect 15349 39149 15458 39152
rect 15401 39097 15458 39149
rect 15349 39094 15458 39097
rect 15349 39091 15401 39094
rect 15458 39088 15516 39094
rect 21352 37832 21410 37838
rect 21467 37832 21519 37835
rect 21410 37829 21519 37832
rect 21410 37777 21467 37829
rect 21410 37774 21519 37777
rect 21352 37768 21410 37774
rect 21467 37771 21519 37774
rect 21767 37829 21819 37835
rect 21767 37771 21819 37777
rect 22067 37829 22119 37835
rect 22067 37771 22119 37777
rect 22367 37829 22419 37835
rect 22367 37771 22419 37777
rect 22667 37829 22719 37835
rect 22667 37771 22719 37777
rect 22967 37829 23019 37835
rect 22967 37771 23019 37777
rect 23267 37829 23319 37835
rect 23267 37771 23319 37777
rect 23567 37829 23619 37835
rect 23858 37832 23916 37838
rect 23567 37771 23619 37777
rect 23776 37774 23858 37832
rect 23858 37768 23916 37774
rect 7722 36791 7780 36797
rect 7780 36733 7892 36791
rect 8049 36788 8101 36794
rect 7722 36727 7780 36733
rect 8049 36730 8101 36736
rect 8349 36788 8401 36794
rect 8349 36730 8401 36736
rect 8649 36788 8701 36794
rect 8649 36730 8701 36736
rect 8949 36788 9001 36794
rect 8949 36730 9001 36736
rect 9249 36788 9301 36794
rect 9249 36730 9301 36736
rect 9549 36788 9601 36794
rect 9549 36730 9601 36736
rect 9849 36788 9901 36794
rect 9849 36730 9901 36736
rect 10149 36791 10201 36794
rect 12922 36791 12980 36797
rect 10149 36788 10278 36791
rect 10201 36736 10278 36788
rect 10149 36733 10278 36736
rect 10336 36733 10342 36791
rect 12980 36733 13092 36791
rect 13249 36788 13301 36794
rect 10149 36730 10201 36733
rect 12922 36727 12980 36733
rect 13249 36730 13301 36736
rect 13549 36788 13601 36794
rect 13549 36730 13601 36736
rect 13849 36788 13901 36794
rect 13849 36730 13901 36736
rect 14149 36788 14201 36794
rect 14149 36730 14201 36736
rect 14449 36788 14501 36794
rect 14449 36730 14501 36736
rect 14749 36788 14801 36794
rect 14749 36730 14801 36736
rect 15049 36788 15101 36794
rect 15049 36730 15101 36736
rect 15349 36791 15401 36794
rect 15349 36788 15478 36791
rect 15401 36736 15478 36788
rect 15349 36733 15478 36736
rect 15536 36733 15542 36791
rect 15349 36730 15401 36733
rect 21326 36706 21396 36712
rect 23882 36706 23952 36712
rect 21396 36642 21492 36700
rect 23776 36642 23882 36700
rect 21326 36630 21396 36636
rect 23882 36630 23952 36636
rect 21346 36496 21416 36502
rect 23853 36496 23923 36502
rect 21416 36432 21492 36490
rect 23776 36432 23853 36490
rect 21346 36420 21416 36426
rect 23853 36420 23923 36426
rect 7752 35659 7810 35665
rect 7810 35601 7892 35659
rect 8063 35656 8115 35662
rect 7752 35595 7810 35601
rect 8063 35598 8115 35604
rect 8363 35656 8415 35662
rect 8363 35598 8415 35604
rect 8663 35656 8715 35662
rect 8663 35598 8715 35604
rect 8963 35656 9015 35662
rect 8963 35598 9015 35604
rect 9263 35656 9315 35662
rect 9263 35598 9315 35604
rect 9563 35656 9615 35662
rect 9563 35598 9615 35604
rect 9863 35656 9915 35662
rect 9863 35598 9915 35604
rect 10163 35659 10215 35662
rect 10258 35659 10316 35665
rect 10163 35656 10258 35659
rect 10215 35604 10258 35656
rect 10163 35601 10258 35604
rect 10163 35598 10215 35601
rect 10258 35595 10316 35601
rect 12952 35659 13010 35665
rect 13010 35601 13092 35659
rect 13263 35656 13315 35662
rect 12952 35595 13010 35601
rect 13263 35598 13315 35604
rect 13563 35656 13615 35662
rect 13563 35598 13615 35604
rect 13863 35656 13915 35662
rect 13863 35598 13915 35604
rect 14163 35656 14215 35662
rect 14163 35598 14215 35604
rect 14463 35656 14515 35662
rect 14463 35598 14515 35604
rect 14763 35656 14815 35662
rect 14763 35598 14815 35604
rect 15063 35656 15115 35662
rect 15063 35598 15115 35604
rect 15363 35659 15415 35662
rect 15458 35659 15516 35665
rect 15363 35656 15458 35659
rect 15415 35604 15458 35656
rect 15363 35601 15458 35604
rect 15363 35598 15415 35601
rect 15458 35595 15516 35601
rect 21332 35358 21390 35364
rect 21466 35358 21518 35361
rect 21390 35355 21518 35358
rect 21390 35303 21466 35355
rect 21390 35300 21518 35303
rect 21332 35294 21390 35300
rect 21466 35297 21518 35300
rect 21766 35355 21818 35361
rect 21766 35297 21818 35303
rect 22066 35355 22118 35361
rect 22066 35297 22118 35303
rect 22366 35355 22418 35361
rect 22366 35297 22418 35303
rect 22666 35355 22718 35361
rect 22666 35297 22718 35303
rect 22966 35355 23018 35361
rect 22966 35297 23018 35303
rect 23266 35355 23318 35361
rect 23266 35297 23318 35303
rect 23566 35355 23618 35361
rect 23888 35358 23946 35364
rect 23566 35297 23618 35303
rect 23776 35300 23888 35358
rect 23888 35294 23946 35300
rect 0 0 200 200
rect 28872 0 29072 200
<< via1 >>
rect 7722 41568 7780 41626
rect 8050 41571 8102 41623
rect 8350 41571 8402 41623
rect 8650 41571 8702 41623
rect 8950 41571 9002 41623
rect 9250 41571 9302 41623
rect 9550 41571 9602 41623
rect 9850 41571 9902 41623
rect 10150 41571 10202 41623
rect 10278 41568 10336 41626
rect 12922 41568 12980 41626
rect 13250 41571 13302 41623
rect 13550 41571 13602 41623
rect 13850 41571 13902 41623
rect 14150 41571 14202 41623
rect 14450 41571 14502 41623
rect 14750 41571 14802 41623
rect 15050 41571 15102 41623
rect 15350 41571 15402 41623
rect 15478 41568 15536 41626
rect 2664 41282 2724 41342
rect 2964 41282 3024 41342
rect 3264 41282 3324 41342
rect 3564 41282 3624 41342
rect 3864 41282 3924 41342
rect 4164 41282 4224 41342
rect 4464 41282 4524 41342
rect 4764 41282 4824 41342
rect 21352 41267 21410 41325
rect 21453 41270 21505 41322
rect 21753 41270 21805 41322
rect 22053 41270 22105 41322
rect 22353 41270 22405 41322
rect 22653 41270 22705 41322
rect 22953 41270 23005 41322
rect 23253 41270 23305 41322
rect 23553 41270 23605 41322
rect 23858 41267 23916 41325
rect 7745 40430 7815 40500
rect 10252 40430 10322 40500
rect 12945 40430 13015 40500
rect 15452 40430 15522 40500
rect 7716 40220 7786 40290
rect 10272 40220 10342 40290
rect 12916 40220 12986 40290
rect 15472 40220 15542 40290
rect 2667 40154 2719 40206
rect 2967 40154 3019 40206
rect 3267 40154 3319 40206
rect 3567 40154 3619 40206
rect 3867 40154 3919 40206
rect 4167 40154 4219 40206
rect 4467 40154 4519 40206
rect 4767 40154 4819 40206
rect 21332 40135 21390 40193
rect 21467 40138 21519 40190
rect 21767 40138 21819 40190
rect 22067 40138 22119 40190
rect 22367 40138 22419 40190
rect 22667 40138 22719 40190
rect 22967 40138 23019 40190
rect 23267 40138 23319 40190
rect 23567 40138 23619 40190
rect 23888 40135 23946 40193
rect 7752 39094 7810 39152
rect 8049 39097 8101 39149
rect 8349 39097 8401 39149
rect 8649 39097 8701 39149
rect 8949 39097 9001 39149
rect 9249 39097 9301 39149
rect 9549 39097 9601 39149
rect 9849 39097 9901 39149
rect 10149 39097 10201 39149
rect 10258 39094 10316 39152
rect 12952 39094 13010 39152
rect 13249 39097 13301 39149
rect 13549 39097 13601 39149
rect 13849 39097 13901 39149
rect 14149 39097 14201 39149
rect 14449 39097 14501 39149
rect 14749 39097 14801 39149
rect 15049 39097 15101 39149
rect 15349 39097 15401 39149
rect 15458 39094 15516 39152
rect 21352 37774 21410 37832
rect 21467 37777 21519 37829
rect 21767 37777 21819 37829
rect 22067 37777 22119 37829
rect 22367 37777 22419 37829
rect 22667 37777 22719 37829
rect 22967 37777 23019 37829
rect 23267 37777 23319 37829
rect 23567 37777 23619 37829
rect 23858 37774 23916 37832
rect 7722 36733 7780 36791
rect 8049 36736 8101 36788
rect 8349 36736 8401 36788
rect 8649 36736 8701 36788
rect 8949 36736 9001 36788
rect 9249 36736 9301 36788
rect 9549 36736 9601 36788
rect 9849 36736 9901 36788
rect 10149 36736 10201 36788
rect 10278 36733 10336 36791
rect 12922 36733 12980 36791
rect 13249 36736 13301 36788
rect 13549 36736 13601 36788
rect 13849 36736 13901 36788
rect 14149 36736 14201 36788
rect 14449 36736 14501 36788
rect 14749 36736 14801 36788
rect 15049 36736 15101 36788
rect 15349 36736 15401 36788
rect 15478 36733 15536 36791
rect 21326 36636 21396 36706
rect 23882 36636 23952 36706
rect 21346 36426 21416 36496
rect 23853 36426 23923 36496
rect 7752 35601 7810 35659
rect 8063 35604 8115 35656
rect 8363 35604 8415 35656
rect 8663 35604 8715 35656
rect 8963 35604 9015 35656
rect 9263 35604 9315 35656
rect 9563 35604 9615 35656
rect 9863 35604 9915 35656
rect 10163 35604 10215 35656
rect 10258 35601 10316 35659
rect 12952 35601 13010 35659
rect 13263 35604 13315 35656
rect 13563 35604 13615 35656
rect 13863 35604 13915 35656
rect 14163 35604 14215 35656
rect 14463 35604 14515 35656
rect 14763 35604 14815 35656
rect 15063 35604 15115 35656
rect 15363 35604 15415 35656
rect 15458 35601 15516 35659
rect 21332 35300 21390 35358
rect 21466 35303 21518 35355
rect 21766 35303 21818 35355
rect 22066 35303 22118 35355
rect 22366 35303 22418 35355
rect 22666 35303 22718 35355
rect 22966 35303 23018 35355
rect 23266 35303 23318 35355
rect 23566 35303 23618 35355
rect 23888 35300 23946 35358
<< metal2 >>
rect 7721 41627 7781 41636
rect 8046 41627 8106 41636
rect 7716 41568 7721 41626
rect 7781 41568 7786 41626
rect 8346 41627 8406 41636
rect 8646 41627 8706 41636
rect 8946 41627 9006 41636
rect 9246 41627 9306 41636
rect 9546 41627 9606 41636
rect 9846 41627 9906 41636
rect 10146 41627 10206 41636
rect 10277 41627 10337 41636
rect 12921 41627 12981 41636
rect 13246 41627 13306 41636
rect 8044 41571 8046 41623
rect 8106 41571 8108 41623
rect 8344 41571 8346 41623
rect 8406 41571 8408 41623
rect 8644 41571 8646 41623
rect 8706 41571 8708 41623
rect 8944 41571 8946 41623
rect 9006 41571 9008 41623
rect 9244 41571 9246 41623
rect 9306 41571 9308 41623
rect 9544 41571 9546 41623
rect 9606 41571 9608 41623
rect 9844 41571 9846 41623
rect 9906 41571 9908 41623
rect 10144 41571 10146 41623
rect 10206 41571 10208 41623
rect 7721 41558 7781 41567
rect 8046 41558 8106 41567
rect 8346 41558 8406 41567
rect 8646 41558 8706 41567
rect 8946 41558 9006 41567
rect 9246 41558 9306 41567
rect 9546 41558 9606 41567
rect 9846 41558 9906 41567
rect 10272 41568 10277 41626
rect 10337 41568 10342 41626
rect 12916 41568 12921 41626
rect 12981 41568 12986 41626
rect 13546 41627 13606 41636
rect 13846 41627 13906 41636
rect 14146 41627 14206 41636
rect 14446 41627 14506 41636
rect 14746 41627 14806 41636
rect 15046 41627 15106 41636
rect 15346 41627 15406 41636
rect 15477 41627 15537 41636
rect 13244 41571 13246 41623
rect 13306 41571 13308 41623
rect 13544 41571 13546 41623
rect 13606 41571 13608 41623
rect 13844 41571 13846 41623
rect 13906 41571 13908 41623
rect 14144 41571 14146 41623
rect 14206 41571 14208 41623
rect 14444 41571 14446 41623
rect 14506 41571 14508 41623
rect 14744 41571 14746 41623
rect 14806 41571 14808 41623
rect 15044 41571 15046 41623
rect 15106 41571 15108 41623
rect 15344 41571 15346 41623
rect 15406 41571 15408 41623
rect 10146 41558 10206 41567
rect 10277 41558 10337 41567
rect 12921 41558 12981 41567
rect 13246 41558 13306 41567
rect 13546 41558 13606 41567
rect 13846 41558 13906 41567
rect 14146 41558 14206 41567
rect 14446 41558 14506 41567
rect 14746 41558 14806 41567
rect 15046 41558 15106 41567
rect 15472 41568 15477 41626
rect 15537 41568 15542 41626
rect 15346 41558 15406 41567
rect 15477 41558 15537 41567
rect 2664 41342 2724 41351
rect 2964 41342 3024 41351
rect 3264 41342 3324 41351
rect 3564 41342 3624 41351
rect 3864 41342 3924 41351
rect 4164 41342 4224 41351
rect 4464 41342 4524 41351
rect 4764 41342 4824 41351
rect 2658 41282 2664 41342
rect 2724 41282 2730 41342
rect 2958 41282 2964 41342
rect 3024 41282 3030 41342
rect 3258 41282 3264 41342
rect 3324 41282 3330 41342
rect 3558 41282 3564 41342
rect 3624 41282 3630 41342
rect 3858 41282 3864 41342
rect 3924 41282 3930 41342
rect 4158 41282 4164 41342
rect 4224 41282 4230 41342
rect 4458 41282 4464 41342
rect 4524 41282 4530 41342
rect 4758 41282 4764 41342
rect 4824 41282 4830 41342
rect 21351 41326 21411 41335
rect 21449 41326 21509 41335
rect 2664 41273 2724 41282
rect 2964 41273 3024 41282
rect 3264 41273 3324 41282
rect 3564 41273 3624 41282
rect 3864 41273 3924 41282
rect 4164 41273 4224 41282
rect 4464 41273 4524 41282
rect 4764 41273 4824 41282
rect 21346 41267 21351 41325
rect 21411 41267 21416 41325
rect 21749 41326 21809 41335
rect 22049 41326 22109 41335
rect 22349 41326 22409 41335
rect 22649 41326 22709 41335
rect 22949 41326 23009 41335
rect 23249 41326 23309 41335
rect 23549 41326 23609 41335
rect 23857 41326 23917 41335
rect 21447 41270 21449 41322
rect 21509 41270 21511 41322
rect 21747 41270 21749 41322
rect 21809 41270 21811 41322
rect 22047 41270 22049 41322
rect 22109 41270 22111 41322
rect 22347 41270 22349 41322
rect 22409 41270 22411 41322
rect 22647 41270 22649 41322
rect 22709 41270 22711 41322
rect 22947 41270 22949 41322
rect 23009 41270 23011 41322
rect 23247 41270 23249 41322
rect 23309 41270 23311 41322
rect 23547 41270 23549 41322
rect 23609 41270 23611 41322
rect 21351 41257 21411 41266
rect 21449 41257 21509 41266
rect 21749 41257 21809 41266
rect 22049 41257 22109 41266
rect 22349 41257 22409 41266
rect 22649 41257 22709 41266
rect 22949 41257 23009 41266
rect 23249 41257 23309 41266
rect 23852 41267 23857 41325
rect 23917 41267 23922 41325
rect 23549 41257 23609 41266
rect 23857 41257 23917 41266
rect 7745 40500 7815 40509
rect 10252 40500 10322 40509
rect 12945 40500 13015 40509
rect 15452 40500 15522 40509
rect 7739 40430 7745 40500
rect 7815 40430 7821 40500
rect 10246 40430 10252 40500
rect 10322 40430 10328 40500
rect 12939 40430 12945 40500
rect 13015 40430 13021 40500
rect 15446 40430 15452 40500
rect 15522 40430 15528 40500
rect 7745 40421 7815 40430
rect 10252 40421 10322 40430
rect 12945 40421 13015 40430
rect 15452 40421 15522 40430
rect 7716 40290 7786 40299
rect 10272 40290 10342 40299
rect 12916 40290 12986 40299
rect 15472 40290 15542 40299
rect 7710 40220 7716 40290
rect 7786 40220 7792 40290
rect 10266 40220 10272 40290
rect 10342 40220 10348 40290
rect 12910 40220 12916 40290
rect 12986 40220 12992 40290
rect 15466 40220 15472 40290
rect 15542 40220 15548 40290
rect 2663 40210 2723 40219
rect 2963 40210 3023 40219
rect 3263 40210 3323 40219
rect 3563 40210 3623 40219
rect 3863 40210 3923 40219
rect 4163 40210 4223 40219
rect 4463 40210 4523 40219
rect 4763 40210 4823 40219
rect 7716 40211 7786 40220
rect 10272 40211 10342 40220
rect 12916 40211 12986 40220
rect 15472 40211 15542 40220
rect 2661 40154 2663 40206
rect 2723 40154 2725 40206
rect 2961 40154 2963 40206
rect 3023 40154 3025 40206
rect 3261 40154 3263 40206
rect 3323 40154 3325 40206
rect 3561 40154 3563 40206
rect 3623 40154 3625 40206
rect 3861 40154 3863 40206
rect 3923 40154 3925 40206
rect 4161 40154 4163 40206
rect 4223 40154 4225 40206
rect 4461 40154 4463 40206
rect 4523 40154 4525 40206
rect 4761 40154 4763 40206
rect 4823 40154 4825 40206
rect 21331 40194 21391 40203
rect 2663 40141 2723 40150
rect 2963 40141 3023 40150
rect 3263 40141 3323 40150
rect 3563 40141 3623 40150
rect 3863 40141 3923 40150
rect 4163 40141 4223 40150
rect 4463 40141 4523 40150
rect 4763 40141 4823 40150
rect 21463 40194 21523 40203
rect 21763 40194 21823 40203
rect 22063 40194 22123 40203
rect 22363 40194 22423 40203
rect 22663 40194 22723 40203
rect 22963 40194 23023 40203
rect 23263 40194 23323 40203
rect 23563 40194 23623 40203
rect 23887 40194 23947 40203
rect 21461 40138 21463 40190
rect 21523 40138 21525 40190
rect 21761 40138 21763 40190
rect 21823 40138 21825 40190
rect 22061 40138 22063 40190
rect 22123 40138 22125 40190
rect 22361 40138 22363 40190
rect 22423 40138 22425 40190
rect 22661 40138 22663 40190
rect 22723 40138 22725 40190
rect 22961 40138 22963 40190
rect 23023 40138 23025 40190
rect 23261 40138 23263 40190
rect 23323 40138 23325 40190
rect 23561 40138 23563 40190
rect 23623 40138 23625 40190
rect 21331 40125 21391 40134
rect 21463 40125 21523 40134
rect 21763 40125 21823 40134
rect 22063 40125 22123 40134
rect 22363 40125 22423 40134
rect 22663 40125 22723 40134
rect 22963 40125 23023 40134
rect 23263 40125 23323 40134
rect 23882 40135 23887 40193
rect 23947 40135 23952 40193
rect 23563 40125 23623 40134
rect 23887 40125 23947 40134
rect 7751 39153 7811 39162
rect 8045 39153 8105 39162
rect 7746 39094 7751 39152
rect 7811 39094 7816 39152
rect 8345 39153 8405 39162
rect 8645 39153 8705 39162
rect 8945 39153 9005 39162
rect 9245 39153 9305 39162
rect 9545 39153 9605 39162
rect 9845 39153 9905 39162
rect 10145 39153 10205 39162
rect 10257 39153 10317 39162
rect 12951 39153 13011 39162
rect 13245 39153 13305 39162
rect 8043 39097 8045 39149
rect 8105 39097 8107 39149
rect 8343 39097 8345 39149
rect 8405 39097 8407 39149
rect 8643 39097 8645 39149
rect 8705 39097 8707 39149
rect 8943 39097 8945 39149
rect 9005 39097 9007 39149
rect 9243 39097 9245 39149
rect 9305 39097 9307 39149
rect 9543 39097 9545 39149
rect 9605 39097 9607 39149
rect 9843 39097 9845 39149
rect 9905 39097 9907 39149
rect 10143 39097 10145 39149
rect 10205 39097 10207 39149
rect 7751 39084 7811 39093
rect 8045 39084 8105 39093
rect 8345 39084 8405 39093
rect 8645 39084 8705 39093
rect 8945 39084 9005 39093
rect 9245 39084 9305 39093
rect 9545 39084 9605 39093
rect 9845 39084 9905 39093
rect 10252 39094 10257 39152
rect 10317 39094 10322 39152
rect 12946 39094 12951 39152
rect 13011 39094 13016 39152
rect 13545 39153 13605 39162
rect 13845 39153 13905 39162
rect 14145 39153 14205 39162
rect 14445 39153 14505 39162
rect 14745 39153 14805 39162
rect 15045 39153 15105 39162
rect 15345 39153 15405 39162
rect 15457 39153 15517 39162
rect 13243 39097 13245 39149
rect 13305 39097 13307 39149
rect 13543 39097 13545 39149
rect 13605 39097 13607 39149
rect 13843 39097 13845 39149
rect 13905 39097 13907 39149
rect 14143 39097 14145 39149
rect 14205 39097 14207 39149
rect 14443 39097 14445 39149
rect 14505 39097 14507 39149
rect 14743 39097 14745 39149
rect 14805 39097 14807 39149
rect 15043 39097 15045 39149
rect 15105 39097 15107 39149
rect 15343 39097 15345 39149
rect 15405 39097 15407 39149
rect 10145 39084 10205 39093
rect 10257 39084 10317 39093
rect 12951 39084 13011 39093
rect 13245 39084 13305 39093
rect 13545 39084 13605 39093
rect 13845 39084 13905 39093
rect 14145 39084 14205 39093
rect 14445 39084 14505 39093
rect 14745 39084 14805 39093
rect 15045 39084 15105 39093
rect 15452 39094 15457 39152
rect 15517 39094 15522 39152
rect 15345 39084 15405 39093
rect 15457 39084 15517 39093
rect 21351 37833 21411 37842
rect 21463 37833 21523 37842
rect 21346 37774 21351 37832
rect 21411 37774 21416 37832
rect 21763 37833 21823 37842
rect 22063 37833 22123 37842
rect 22363 37833 22423 37842
rect 22663 37833 22723 37842
rect 22963 37833 23023 37842
rect 23263 37833 23323 37842
rect 23563 37833 23623 37842
rect 23857 37833 23917 37842
rect 21461 37777 21463 37829
rect 21523 37777 21525 37829
rect 21761 37777 21763 37829
rect 21823 37777 21825 37829
rect 22061 37777 22063 37829
rect 22123 37777 22125 37829
rect 22361 37777 22363 37829
rect 22423 37777 22425 37829
rect 22661 37777 22663 37829
rect 22723 37777 22725 37829
rect 22961 37777 22963 37829
rect 23023 37777 23025 37829
rect 23261 37777 23263 37829
rect 23323 37777 23325 37829
rect 23561 37777 23563 37829
rect 23623 37777 23625 37829
rect 21351 37764 21411 37773
rect 21463 37764 21523 37773
rect 21763 37764 21823 37773
rect 22063 37764 22123 37773
rect 22363 37764 22423 37773
rect 22663 37764 22723 37773
rect 22963 37764 23023 37773
rect 23263 37764 23323 37773
rect 23852 37774 23857 37832
rect 23917 37774 23922 37832
rect 23563 37764 23623 37773
rect 23857 37764 23917 37773
rect 7721 36792 7781 36801
rect 8045 36792 8105 36801
rect 7716 36733 7721 36791
rect 7781 36733 7786 36791
rect 8345 36792 8405 36801
rect 8645 36792 8705 36801
rect 8945 36792 9005 36801
rect 9245 36792 9305 36801
rect 9545 36792 9605 36801
rect 9845 36792 9905 36801
rect 10145 36792 10205 36801
rect 10277 36792 10337 36801
rect 12921 36792 12981 36801
rect 13245 36792 13305 36801
rect 8043 36736 8045 36788
rect 8105 36736 8107 36788
rect 8343 36736 8345 36788
rect 8405 36736 8407 36788
rect 8643 36736 8645 36788
rect 8705 36736 8707 36788
rect 8943 36736 8945 36788
rect 9005 36736 9007 36788
rect 9243 36736 9245 36788
rect 9305 36736 9307 36788
rect 9543 36736 9545 36788
rect 9605 36736 9607 36788
rect 9843 36736 9845 36788
rect 9905 36736 9907 36788
rect 10143 36736 10145 36788
rect 10205 36736 10207 36788
rect 7721 36723 7781 36732
rect 8045 36723 8105 36732
rect 8345 36723 8405 36732
rect 8645 36723 8705 36732
rect 8945 36723 9005 36732
rect 9245 36723 9305 36732
rect 9545 36723 9605 36732
rect 9845 36723 9905 36732
rect 10145 36723 10205 36732
rect 12916 36733 12921 36791
rect 12981 36733 12986 36791
rect 13545 36792 13605 36801
rect 13845 36792 13905 36801
rect 14145 36792 14205 36801
rect 14445 36792 14505 36801
rect 14745 36792 14805 36801
rect 15045 36792 15105 36801
rect 15345 36792 15405 36801
rect 15477 36792 15537 36801
rect 13243 36736 13245 36788
rect 13305 36736 13307 36788
rect 13543 36736 13545 36788
rect 13605 36736 13607 36788
rect 13843 36736 13845 36788
rect 13905 36736 13907 36788
rect 14143 36736 14145 36788
rect 14205 36736 14207 36788
rect 14443 36736 14445 36788
rect 14505 36736 14507 36788
rect 14743 36736 14745 36788
rect 14805 36736 14807 36788
rect 15043 36736 15045 36788
rect 15105 36736 15107 36788
rect 15343 36736 15345 36788
rect 15405 36736 15407 36788
rect 10277 36723 10337 36732
rect 12921 36723 12981 36732
rect 13245 36723 13305 36732
rect 13545 36723 13605 36732
rect 13845 36723 13905 36732
rect 14145 36723 14205 36732
rect 14445 36723 14505 36732
rect 14745 36723 14805 36732
rect 15045 36723 15105 36732
rect 15345 36723 15405 36732
rect 15477 36723 15537 36732
rect 21326 36706 21396 36715
rect 23882 36706 23952 36715
rect 21320 36636 21326 36706
rect 21396 36636 21402 36706
rect 23876 36636 23882 36706
rect 23952 36636 23958 36706
rect 21326 36627 21396 36636
rect 23882 36627 23952 36636
rect 21346 36496 21416 36505
rect 23853 36496 23923 36505
rect 21340 36426 21346 36496
rect 21416 36426 21422 36496
rect 23847 36426 23853 36496
rect 23923 36426 23929 36496
rect 21346 36417 21416 36426
rect 23853 36417 23923 36426
rect 7751 35660 7811 35669
rect 8059 35660 8119 35669
rect 7746 35601 7751 35659
rect 7811 35601 7816 35659
rect 8359 35660 8419 35669
rect 8659 35660 8719 35669
rect 8959 35660 9019 35669
rect 9259 35660 9319 35669
rect 9559 35660 9619 35669
rect 9859 35660 9919 35669
rect 10159 35660 10219 35669
rect 10257 35660 10317 35669
rect 12951 35660 13011 35669
rect 13259 35660 13319 35669
rect 8057 35604 8059 35656
rect 8119 35604 8121 35656
rect 8357 35604 8359 35656
rect 8419 35604 8421 35656
rect 8657 35604 8659 35656
rect 8719 35604 8721 35656
rect 8957 35604 8959 35656
rect 9019 35604 9021 35656
rect 9257 35604 9259 35656
rect 9319 35604 9321 35656
rect 9557 35604 9559 35656
rect 9619 35604 9621 35656
rect 9857 35604 9859 35656
rect 9919 35604 9921 35656
rect 10157 35604 10159 35656
rect 10219 35604 10221 35656
rect 7751 35591 7811 35600
rect 8059 35591 8119 35600
rect 8359 35591 8419 35600
rect 8659 35591 8719 35600
rect 8959 35591 9019 35600
rect 9259 35591 9319 35600
rect 9559 35591 9619 35600
rect 9859 35591 9919 35600
rect 10252 35601 10257 35659
rect 10317 35601 10322 35659
rect 12946 35601 12951 35659
rect 13011 35601 13016 35659
rect 13559 35660 13619 35669
rect 13859 35660 13919 35669
rect 14159 35660 14219 35669
rect 14459 35660 14519 35669
rect 14759 35660 14819 35669
rect 15059 35660 15119 35669
rect 15359 35660 15419 35669
rect 15457 35660 15517 35669
rect 13257 35604 13259 35656
rect 13319 35604 13321 35656
rect 13557 35604 13559 35656
rect 13619 35604 13621 35656
rect 13857 35604 13859 35656
rect 13919 35604 13921 35656
rect 14157 35604 14159 35656
rect 14219 35604 14221 35656
rect 14457 35604 14459 35656
rect 14519 35604 14521 35656
rect 14757 35604 14759 35656
rect 14819 35604 14821 35656
rect 15057 35604 15059 35656
rect 15119 35604 15121 35656
rect 15357 35604 15359 35656
rect 15419 35604 15421 35656
rect 10159 35591 10219 35600
rect 10257 35591 10317 35600
rect 12951 35591 13011 35600
rect 13259 35591 13319 35600
rect 13559 35591 13619 35600
rect 13859 35591 13919 35600
rect 14159 35591 14219 35600
rect 14459 35591 14519 35600
rect 14759 35591 14819 35600
rect 15059 35591 15119 35600
rect 15452 35601 15457 35659
rect 15517 35601 15522 35659
rect 15359 35591 15419 35600
rect 15457 35591 15517 35600
rect 21331 35359 21391 35368
rect 21462 35359 21522 35368
rect 21326 35300 21331 35358
rect 21391 35300 21396 35358
rect 21762 35359 21822 35368
rect 22062 35359 22122 35368
rect 22362 35359 22422 35368
rect 22662 35359 22722 35368
rect 22962 35359 23022 35368
rect 23262 35359 23322 35368
rect 23562 35359 23622 35368
rect 23887 35359 23947 35368
rect 21460 35303 21462 35355
rect 21522 35303 21524 35355
rect 21760 35303 21762 35355
rect 21822 35303 21824 35355
rect 22060 35303 22062 35355
rect 22122 35303 22124 35355
rect 22360 35303 22362 35355
rect 22422 35303 22424 35355
rect 22660 35303 22662 35355
rect 22722 35303 22724 35355
rect 22960 35303 22962 35355
rect 23022 35303 23024 35355
rect 23260 35303 23262 35355
rect 23322 35303 23324 35355
rect 23560 35303 23562 35355
rect 23622 35303 23624 35355
rect 21331 35290 21391 35299
rect 21462 35290 21522 35299
rect 21762 35290 21822 35299
rect 22062 35290 22122 35299
rect 22362 35290 22422 35299
rect 22662 35290 22722 35299
rect 22962 35290 23022 35299
rect 23262 35290 23322 35299
rect 23882 35300 23887 35358
rect 23947 35300 23952 35358
rect 23562 35290 23622 35299
rect 23887 35290 23947 35299
rect 13131 19974 13269 19983
rect 13131 19074 13269 19836
rect 14131 17388 14269 17397
rect 13693 17250 14131 17388
rect 14131 17241 14269 17250
rect 13131 10969 13269 10978
rect 13131 9734 13269 10831
rect 13684 7843 13693 7981
rect 13831 7843 13840 7981
rect 17354 6419 17492 6428
rect 17354 6272 17492 6281
rect 17354 4595 17492 4604
rect 17354 4448 17492 4457
<< via2 >>
rect 7721 41626 7781 41627
rect 7721 41568 7722 41626
rect 7722 41568 7780 41626
rect 7780 41568 7781 41626
rect 8046 41623 8106 41627
rect 8346 41623 8406 41627
rect 8646 41623 8706 41627
rect 8946 41623 9006 41627
rect 9246 41623 9306 41627
rect 9546 41623 9606 41627
rect 9846 41623 9906 41627
rect 10146 41623 10206 41627
rect 10277 41626 10337 41627
rect 12921 41626 12981 41627
rect 8046 41571 8050 41623
rect 8050 41571 8102 41623
rect 8102 41571 8106 41623
rect 8346 41571 8350 41623
rect 8350 41571 8402 41623
rect 8402 41571 8406 41623
rect 8646 41571 8650 41623
rect 8650 41571 8702 41623
rect 8702 41571 8706 41623
rect 8946 41571 8950 41623
rect 8950 41571 9002 41623
rect 9002 41571 9006 41623
rect 9246 41571 9250 41623
rect 9250 41571 9302 41623
rect 9302 41571 9306 41623
rect 9546 41571 9550 41623
rect 9550 41571 9602 41623
rect 9602 41571 9606 41623
rect 9846 41571 9850 41623
rect 9850 41571 9902 41623
rect 9902 41571 9906 41623
rect 10146 41571 10150 41623
rect 10150 41571 10202 41623
rect 10202 41571 10206 41623
rect 7721 41567 7781 41568
rect 8046 41567 8106 41571
rect 8346 41567 8406 41571
rect 8646 41567 8706 41571
rect 8946 41567 9006 41571
rect 9246 41567 9306 41571
rect 9546 41567 9606 41571
rect 9846 41567 9906 41571
rect 10146 41567 10206 41571
rect 10277 41568 10278 41626
rect 10278 41568 10336 41626
rect 10336 41568 10337 41626
rect 12921 41568 12922 41626
rect 12922 41568 12980 41626
rect 12980 41568 12981 41626
rect 13246 41623 13306 41627
rect 13546 41623 13606 41627
rect 13846 41623 13906 41627
rect 14146 41623 14206 41627
rect 14446 41623 14506 41627
rect 14746 41623 14806 41627
rect 15046 41623 15106 41627
rect 15346 41623 15406 41627
rect 15477 41626 15537 41627
rect 13246 41571 13250 41623
rect 13250 41571 13302 41623
rect 13302 41571 13306 41623
rect 13546 41571 13550 41623
rect 13550 41571 13602 41623
rect 13602 41571 13606 41623
rect 13846 41571 13850 41623
rect 13850 41571 13902 41623
rect 13902 41571 13906 41623
rect 14146 41571 14150 41623
rect 14150 41571 14202 41623
rect 14202 41571 14206 41623
rect 14446 41571 14450 41623
rect 14450 41571 14502 41623
rect 14502 41571 14506 41623
rect 14746 41571 14750 41623
rect 14750 41571 14802 41623
rect 14802 41571 14806 41623
rect 15046 41571 15050 41623
rect 15050 41571 15102 41623
rect 15102 41571 15106 41623
rect 15346 41571 15350 41623
rect 15350 41571 15402 41623
rect 15402 41571 15406 41623
rect 10277 41567 10337 41568
rect 12921 41567 12981 41568
rect 13246 41567 13306 41571
rect 13546 41567 13606 41571
rect 13846 41567 13906 41571
rect 14146 41567 14206 41571
rect 14446 41567 14506 41571
rect 14746 41567 14806 41571
rect 15046 41567 15106 41571
rect 15346 41567 15406 41571
rect 15477 41568 15478 41626
rect 15478 41568 15536 41626
rect 15536 41568 15537 41626
rect 15477 41567 15537 41568
rect 2664 41282 2724 41342
rect 2964 41282 3024 41342
rect 3264 41282 3324 41342
rect 3564 41282 3624 41342
rect 3864 41282 3924 41342
rect 4164 41282 4224 41342
rect 4464 41282 4524 41342
rect 4764 41282 4824 41342
rect 21351 41325 21411 41326
rect 21351 41267 21352 41325
rect 21352 41267 21410 41325
rect 21410 41267 21411 41325
rect 21449 41322 21509 41326
rect 21749 41322 21809 41326
rect 22049 41322 22109 41326
rect 22349 41322 22409 41326
rect 22649 41322 22709 41326
rect 22949 41322 23009 41326
rect 23249 41322 23309 41326
rect 23549 41322 23609 41326
rect 23857 41325 23917 41326
rect 21449 41270 21453 41322
rect 21453 41270 21505 41322
rect 21505 41270 21509 41322
rect 21749 41270 21753 41322
rect 21753 41270 21805 41322
rect 21805 41270 21809 41322
rect 22049 41270 22053 41322
rect 22053 41270 22105 41322
rect 22105 41270 22109 41322
rect 22349 41270 22353 41322
rect 22353 41270 22405 41322
rect 22405 41270 22409 41322
rect 22649 41270 22653 41322
rect 22653 41270 22705 41322
rect 22705 41270 22709 41322
rect 22949 41270 22953 41322
rect 22953 41270 23005 41322
rect 23005 41270 23009 41322
rect 23249 41270 23253 41322
rect 23253 41270 23305 41322
rect 23305 41270 23309 41322
rect 23549 41270 23553 41322
rect 23553 41270 23605 41322
rect 23605 41270 23609 41322
rect 21351 41266 21411 41267
rect 21449 41266 21509 41270
rect 21749 41266 21809 41270
rect 22049 41266 22109 41270
rect 22349 41266 22409 41270
rect 22649 41266 22709 41270
rect 22949 41266 23009 41270
rect 23249 41266 23309 41270
rect 23549 41266 23609 41270
rect 23857 41267 23858 41325
rect 23858 41267 23916 41325
rect 23916 41267 23917 41325
rect 23857 41266 23917 41267
rect 7745 40430 7815 40500
rect 10252 40430 10322 40500
rect 12945 40430 13015 40500
rect 15452 40430 15522 40500
rect 7716 40220 7786 40290
rect 10272 40220 10342 40290
rect 12916 40220 12986 40290
rect 15472 40220 15542 40290
rect 2663 40206 2723 40210
rect 2963 40206 3023 40210
rect 3263 40206 3323 40210
rect 3563 40206 3623 40210
rect 3863 40206 3923 40210
rect 4163 40206 4223 40210
rect 4463 40206 4523 40210
rect 4763 40206 4823 40210
rect 2663 40154 2667 40206
rect 2667 40154 2719 40206
rect 2719 40154 2723 40206
rect 2963 40154 2967 40206
rect 2967 40154 3019 40206
rect 3019 40154 3023 40206
rect 3263 40154 3267 40206
rect 3267 40154 3319 40206
rect 3319 40154 3323 40206
rect 3563 40154 3567 40206
rect 3567 40154 3619 40206
rect 3619 40154 3623 40206
rect 3863 40154 3867 40206
rect 3867 40154 3919 40206
rect 3919 40154 3923 40206
rect 4163 40154 4167 40206
rect 4167 40154 4219 40206
rect 4219 40154 4223 40206
rect 4463 40154 4467 40206
rect 4467 40154 4519 40206
rect 4519 40154 4523 40206
rect 4763 40154 4767 40206
rect 4767 40154 4819 40206
rect 4819 40154 4823 40206
rect 21331 40193 21391 40194
rect 2663 40150 2723 40154
rect 2963 40150 3023 40154
rect 3263 40150 3323 40154
rect 3563 40150 3623 40154
rect 3863 40150 3923 40154
rect 4163 40150 4223 40154
rect 4463 40150 4523 40154
rect 4763 40150 4823 40154
rect 21331 40135 21332 40193
rect 21332 40135 21390 40193
rect 21390 40135 21391 40193
rect 21463 40190 21523 40194
rect 21763 40190 21823 40194
rect 22063 40190 22123 40194
rect 22363 40190 22423 40194
rect 22663 40190 22723 40194
rect 22963 40190 23023 40194
rect 23263 40190 23323 40194
rect 23563 40190 23623 40194
rect 23887 40193 23947 40194
rect 21463 40138 21467 40190
rect 21467 40138 21519 40190
rect 21519 40138 21523 40190
rect 21763 40138 21767 40190
rect 21767 40138 21819 40190
rect 21819 40138 21823 40190
rect 22063 40138 22067 40190
rect 22067 40138 22119 40190
rect 22119 40138 22123 40190
rect 22363 40138 22367 40190
rect 22367 40138 22419 40190
rect 22419 40138 22423 40190
rect 22663 40138 22667 40190
rect 22667 40138 22719 40190
rect 22719 40138 22723 40190
rect 22963 40138 22967 40190
rect 22967 40138 23019 40190
rect 23019 40138 23023 40190
rect 23263 40138 23267 40190
rect 23267 40138 23319 40190
rect 23319 40138 23323 40190
rect 23563 40138 23567 40190
rect 23567 40138 23619 40190
rect 23619 40138 23623 40190
rect 21331 40134 21391 40135
rect 21463 40134 21523 40138
rect 21763 40134 21823 40138
rect 22063 40134 22123 40138
rect 22363 40134 22423 40138
rect 22663 40134 22723 40138
rect 22963 40134 23023 40138
rect 23263 40134 23323 40138
rect 23563 40134 23623 40138
rect 23887 40135 23888 40193
rect 23888 40135 23946 40193
rect 23946 40135 23947 40193
rect 23887 40134 23947 40135
rect 7751 39152 7811 39153
rect 7751 39094 7752 39152
rect 7752 39094 7810 39152
rect 7810 39094 7811 39152
rect 8045 39149 8105 39153
rect 8345 39149 8405 39153
rect 8645 39149 8705 39153
rect 8945 39149 9005 39153
rect 9245 39149 9305 39153
rect 9545 39149 9605 39153
rect 9845 39149 9905 39153
rect 10145 39149 10205 39153
rect 10257 39152 10317 39153
rect 12951 39152 13011 39153
rect 8045 39097 8049 39149
rect 8049 39097 8101 39149
rect 8101 39097 8105 39149
rect 8345 39097 8349 39149
rect 8349 39097 8401 39149
rect 8401 39097 8405 39149
rect 8645 39097 8649 39149
rect 8649 39097 8701 39149
rect 8701 39097 8705 39149
rect 8945 39097 8949 39149
rect 8949 39097 9001 39149
rect 9001 39097 9005 39149
rect 9245 39097 9249 39149
rect 9249 39097 9301 39149
rect 9301 39097 9305 39149
rect 9545 39097 9549 39149
rect 9549 39097 9601 39149
rect 9601 39097 9605 39149
rect 9845 39097 9849 39149
rect 9849 39097 9901 39149
rect 9901 39097 9905 39149
rect 10145 39097 10149 39149
rect 10149 39097 10201 39149
rect 10201 39097 10205 39149
rect 7751 39093 7811 39094
rect 8045 39093 8105 39097
rect 8345 39093 8405 39097
rect 8645 39093 8705 39097
rect 8945 39093 9005 39097
rect 9245 39093 9305 39097
rect 9545 39093 9605 39097
rect 9845 39093 9905 39097
rect 10145 39093 10205 39097
rect 10257 39094 10258 39152
rect 10258 39094 10316 39152
rect 10316 39094 10317 39152
rect 12951 39094 12952 39152
rect 12952 39094 13010 39152
rect 13010 39094 13011 39152
rect 13245 39149 13305 39153
rect 13545 39149 13605 39153
rect 13845 39149 13905 39153
rect 14145 39149 14205 39153
rect 14445 39149 14505 39153
rect 14745 39149 14805 39153
rect 15045 39149 15105 39153
rect 15345 39149 15405 39153
rect 15457 39152 15517 39153
rect 13245 39097 13249 39149
rect 13249 39097 13301 39149
rect 13301 39097 13305 39149
rect 13545 39097 13549 39149
rect 13549 39097 13601 39149
rect 13601 39097 13605 39149
rect 13845 39097 13849 39149
rect 13849 39097 13901 39149
rect 13901 39097 13905 39149
rect 14145 39097 14149 39149
rect 14149 39097 14201 39149
rect 14201 39097 14205 39149
rect 14445 39097 14449 39149
rect 14449 39097 14501 39149
rect 14501 39097 14505 39149
rect 14745 39097 14749 39149
rect 14749 39097 14801 39149
rect 14801 39097 14805 39149
rect 15045 39097 15049 39149
rect 15049 39097 15101 39149
rect 15101 39097 15105 39149
rect 15345 39097 15349 39149
rect 15349 39097 15401 39149
rect 15401 39097 15405 39149
rect 10257 39093 10317 39094
rect 12951 39093 13011 39094
rect 13245 39093 13305 39097
rect 13545 39093 13605 39097
rect 13845 39093 13905 39097
rect 14145 39093 14205 39097
rect 14445 39093 14505 39097
rect 14745 39093 14805 39097
rect 15045 39093 15105 39097
rect 15345 39093 15405 39097
rect 15457 39094 15458 39152
rect 15458 39094 15516 39152
rect 15516 39094 15517 39152
rect 15457 39093 15517 39094
rect 21351 37832 21411 37833
rect 21351 37774 21352 37832
rect 21352 37774 21410 37832
rect 21410 37774 21411 37832
rect 21463 37829 21523 37833
rect 21763 37829 21823 37833
rect 22063 37829 22123 37833
rect 22363 37829 22423 37833
rect 22663 37829 22723 37833
rect 22963 37829 23023 37833
rect 23263 37829 23323 37833
rect 23563 37829 23623 37833
rect 23857 37832 23917 37833
rect 21463 37777 21467 37829
rect 21467 37777 21519 37829
rect 21519 37777 21523 37829
rect 21763 37777 21767 37829
rect 21767 37777 21819 37829
rect 21819 37777 21823 37829
rect 22063 37777 22067 37829
rect 22067 37777 22119 37829
rect 22119 37777 22123 37829
rect 22363 37777 22367 37829
rect 22367 37777 22419 37829
rect 22419 37777 22423 37829
rect 22663 37777 22667 37829
rect 22667 37777 22719 37829
rect 22719 37777 22723 37829
rect 22963 37777 22967 37829
rect 22967 37777 23019 37829
rect 23019 37777 23023 37829
rect 23263 37777 23267 37829
rect 23267 37777 23319 37829
rect 23319 37777 23323 37829
rect 23563 37777 23567 37829
rect 23567 37777 23619 37829
rect 23619 37777 23623 37829
rect 21351 37773 21411 37774
rect 21463 37773 21523 37777
rect 21763 37773 21823 37777
rect 22063 37773 22123 37777
rect 22363 37773 22423 37777
rect 22663 37773 22723 37777
rect 22963 37773 23023 37777
rect 23263 37773 23323 37777
rect 23563 37773 23623 37777
rect 23857 37774 23858 37832
rect 23858 37774 23916 37832
rect 23916 37774 23917 37832
rect 23857 37773 23917 37774
rect 7721 36791 7781 36792
rect 7721 36733 7722 36791
rect 7722 36733 7780 36791
rect 7780 36733 7781 36791
rect 8045 36788 8105 36792
rect 8345 36788 8405 36792
rect 8645 36788 8705 36792
rect 8945 36788 9005 36792
rect 9245 36788 9305 36792
rect 9545 36788 9605 36792
rect 9845 36788 9905 36792
rect 10145 36788 10205 36792
rect 10277 36791 10337 36792
rect 12921 36791 12981 36792
rect 8045 36736 8049 36788
rect 8049 36736 8101 36788
rect 8101 36736 8105 36788
rect 8345 36736 8349 36788
rect 8349 36736 8401 36788
rect 8401 36736 8405 36788
rect 8645 36736 8649 36788
rect 8649 36736 8701 36788
rect 8701 36736 8705 36788
rect 8945 36736 8949 36788
rect 8949 36736 9001 36788
rect 9001 36736 9005 36788
rect 9245 36736 9249 36788
rect 9249 36736 9301 36788
rect 9301 36736 9305 36788
rect 9545 36736 9549 36788
rect 9549 36736 9601 36788
rect 9601 36736 9605 36788
rect 9845 36736 9849 36788
rect 9849 36736 9901 36788
rect 9901 36736 9905 36788
rect 10145 36736 10149 36788
rect 10149 36736 10201 36788
rect 10201 36736 10205 36788
rect 7721 36732 7781 36733
rect 8045 36732 8105 36736
rect 8345 36732 8405 36736
rect 8645 36732 8705 36736
rect 8945 36732 9005 36736
rect 9245 36732 9305 36736
rect 9545 36732 9605 36736
rect 9845 36732 9905 36736
rect 10145 36732 10205 36736
rect 10277 36733 10278 36791
rect 10278 36733 10336 36791
rect 10336 36733 10337 36791
rect 12921 36733 12922 36791
rect 12922 36733 12980 36791
rect 12980 36733 12981 36791
rect 13245 36788 13305 36792
rect 13545 36788 13605 36792
rect 13845 36788 13905 36792
rect 14145 36788 14205 36792
rect 14445 36788 14505 36792
rect 14745 36788 14805 36792
rect 15045 36788 15105 36792
rect 15345 36788 15405 36792
rect 15477 36791 15537 36792
rect 13245 36736 13249 36788
rect 13249 36736 13301 36788
rect 13301 36736 13305 36788
rect 13545 36736 13549 36788
rect 13549 36736 13601 36788
rect 13601 36736 13605 36788
rect 13845 36736 13849 36788
rect 13849 36736 13901 36788
rect 13901 36736 13905 36788
rect 14145 36736 14149 36788
rect 14149 36736 14201 36788
rect 14201 36736 14205 36788
rect 14445 36736 14449 36788
rect 14449 36736 14501 36788
rect 14501 36736 14505 36788
rect 14745 36736 14749 36788
rect 14749 36736 14801 36788
rect 14801 36736 14805 36788
rect 15045 36736 15049 36788
rect 15049 36736 15101 36788
rect 15101 36736 15105 36788
rect 15345 36736 15349 36788
rect 15349 36736 15401 36788
rect 15401 36736 15405 36788
rect 10277 36732 10337 36733
rect 12921 36732 12981 36733
rect 13245 36732 13305 36736
rect 13545 36732 13605 36736
rect 13845 36732 13905 36736
rect 14145 36732 14205 36736
rect 14445 36732 14505 36736
rect 14745 36732 14805 36736
rect 15045 36732 15105 36736
rect 15345 36732 15405 36736
rect 15477 36733 15478 36791
rect 15478 36733 15536 36791
rect 15536 36733 15537 36791
rect 15477 36732 15537 36733
rect 21326 36636 21396 36706
rect 23882 36636 23952 36706
rect 21346 36426 21416 36496
rect 23853 36426 23923 36496
rect 7751 35659 7811 35660
rect 7751 35601 7752 35659
rect 7752 35601 7810 35659
rect 7810 35601 7811 35659
rect 8059 35656 8119 35660
rect 8359 35656 8419 35660
rect 8659 35656 8719 35660
rect 8959 35656 9019 35660
rect 9259 35656 9319 35660
rect 9559 35656 9619 35660
rect 9859 35656 9919 35660
rect 10159 35656 10219 35660
rect 10257 35659 10317 35660
rect 12951 35659 13011 35660
rect 8059 35604 8063 35656
rect 8063 35604 8115 35656
rect 8115 35604 8119 35656
rect 8359 35604 8363 35656
rect 8363 35604 8415 35656
rect 8415 35604 8419 35656
rect 8659 35604 8663 35656
rect 8663 35604 8715 35656
rect 8715 35604 8719 35656
rect 8959 35604 8963 35656
rect 8963 35604 9015 35656
rect 9015 35604 9019 35656
rect 9259 35604 9263 35656
rect 9263 35604 9315 35656
rect 9315 35604 9319 35656
rect 9559 35604 9563 35656
rect 9563 35604 9615 35656
rect 9615 35604 9619 35656
rect 9859 35604 9863 35656
rect 9863 35604 9915 35656
rect 9915 35604 9919 35656
rect 10159 35604 10163 35656
rect 10163 35604 10215 35656
rect 10215 35604 10219 35656
rect 7751 35600 7811 35601
rect 8059 35600 8119 35604
rect 8359 35600 8419 35604
rect 8659 35600 8719 35604
rect 8959 35600 9019 35604
rect 9259 35600 9319 35604
rect 9559 35600 9619 35604
rect 9859 35600 9919 35604
rect 10159 35600 10219 35604
rect 10257 35601 10258 35659
rect 10258 35601 10316 35659
rect 10316 35601 10317 35659
rect 12951 35601 12952 35659
rect 12952 35601 13010 35659
rect 13010 35601 13011 35659
rect 13259 35656 13319 35660
rect 13559 35656 13619 35660
rect 13859 35656 13919 35660
rect 14159 35656 14219 35660
rect 14459 35656 14519 35660
rect 14759 35656 14819 35660
rect 15059 35656 15119 35660
rect 15359 35656 15419 35660
rect 15457 35659 15517 35660
rect 13259 35604 13263 35656
rect 13263 35604 13315 35656
rect 13315 35604 13319 35656
rect 13559 35604 13563 35656
rect 13563 35604 13615 35656
rect 13615 35604 13619 35656
rect 13859 35604 13863 35656
rect 13863 35604 13915 35656
rect 13915 35604 13919 35656
rect 14159 35604 14163 35656
rect 14163 35604 14215 35656
rect 14215 35604 14219 35656
rect 14459 35604 14463 35656
rect 14463 35604 14515 35656
rect 14515 35604 14519 35656
rect 14759 35604 14763 35656
rect 14763 35604 14815 35656
rect 14815 35604 14819 35656
rect 15059 35604 15063 35656
rect 15063 35604 15115 35656
rect 15115 35604 15119 35656
rect 15359 35604 15363 35656
rect 15363 35604 15415 35656
rect 15415 35604 15419 35656
rect 10257 35600 10317 35601
rect 12951 35600 13011 35601
rect 13259 35600 13319 35604
rect 13559 35600 13619 35604
rect 13859 35600 13919 35604
rect 14159 35600 14219 35604
rect 14459 35600 14519 35604
rect 14759 35600 14819 35604
rect 15059 35600 15119 35604
rect 15359 35600 15419 35604
rect 15457 35601 15458 35659
rect 15458 35601 15516 35659
rect 15516 35601 15517 35659
rect 15457 35600 15517 35601
rect 21331 35358 21391 35359
rect 21331 35300 21332 35358
rect 21332 35300 21390 35358
rect 21390 35300 21391 35358
rect 21462 35355 21522 35359
rect 21762 35355 21822 35359
rect 22062 35355 22122 35359
rect 22362 35355 22422 35359
rect 22662 35355 22722 35359
rect 22962 35355 23022 35359
rect 23262 35355 23322 35359
rect 23562 35355 23622 35359
rect 23887 35358 23947 35359
rect 21462 35303 21466 35355
rect 21466 35303 21518 35355
rect 21518 35303 21522 35355
rect 21762 35303 21766 35355
rect 21766 35303 21818 35355
rect 21818 35303 21822 35355
rect 22062 35303 22066 35355
rect 22066 35303 22118 35355
rect 22118 35303 22122 35355
rect 22362 35303 22366 35355
rect 22366 35303 22418 35355
rect 22418 35303 22422 35355
rect 22662 35303 22666 35355
rect 22666 35303 22718 35355
rect 22718 35303 22722 35355
rect 22962 35303 22966 35355
rect 22966 35303 23018 35355
rect 23018 35303 23022 35355
rect 23262 35303 23266 35355
rect 23266 35303 23318 35355
rect 23318 35303 23322 35355
rect 23562 35303 23566 35355
rect 23566 35303 23618 35355
rect 23618 35303 23622 35355
rect 21331 35299 21391 35300
rect 21462 35299 21522 35303
rect 21762 35299 21822 35303
rect 22062 35299 22122 35303
rect 22362 35299 22422 35303
rect 22662 35299 22722 35303
rect 22962 35299 23022 35303
rect 23262 35299 23322 35303
rect 23562 35299 23622 35303
rect 23887 35300 23888 35358
rect 23888 35300 23946 35358
rect 23946 35300 23947 35358
rect 23887 35299 23947 35300
rect 13131 19836 13269 19974
rect 14131 17250 14269 17388
rect 13131 10831 13269 10969
rect 13693 7843 13831 7981
rect 17354 6281 17492 6419
rect 17354 4457 17492 4595
<< metal3 >>
rect 7800 41637 8200 41638
rect 8800 41637 9200 41638
rect 9800 41637 10200 41638
rect 13000 41637 13400 41638
rect 14000 41637 14400 41638
rect 15000 41637 15400 41638
rect 7711 41632 10347 41637
rect 7711 41627 8800 41632
rect 9200 41627 10347 41632
rect 7711 41567 7721 41627
rect 7781 41567 8046 41627
rect 8106 41567 8346 41627
rect 8406 41567 8646 41627
rect 8706 41567 8800 41627
rect 9200 41567 9246 41627
rect 9306 41567 9546 41627
rect 9606 41567 9846 41627
rect 9906 41567 10146 41627
rect 10206 41567 10277 41627
rect 10337 41567 10347 41627
rect 7711 41562 8800 41567
rect 9200 41562 10347 41567
rect 7711 41557 10347 41562
rect 12911 41632 15547 41637
rect 12911 41627 14000 41632
rect 14400 41627 15547 41632
rect 12911 41567 12921 41627
rect 12981 41567 13246 41627
rect 13306 41567 13546 41627
rect 13606 41567 13846 41627
rect 13906 41567 14000 41627
rect 14400 41567 14446 41627
rect 14506 41567 14746 41627
rect 14806 41567 15046 41627
rect 15106 41567 15346 41627
rect 15406 41567 15477 41627
rect 15537 41567 15547 41627
rect 12911 41562 14000 41567
rect 14400 41562 15547 41567
rect 12911 41557 15547 41562
rect 7800 41556 8200 41557
rect 8800 41556 9200 41557
rect 9800 41556 10200 41557
rect 13000 41556 13400 41557
rect 14000 41556 14400 41557
rect 15000 41556 15400 41557
rect 4200 41347 4600 41353
rect 2659 41342 4200 41347
rect 4600 41342 4829 41347
rect 2659 41282 2664 41342
rect 2724 41282 2964 41342
rect 3024 41282 3264 41342
rect 3324 41282 3564 41342
rect 3624 41282 3864 41342
rect 3924 41282 4164 41342
rect 4600 41282 4764 41342
rect 4824 41282 4829 41342
rect 21400 41331 21800 41337
rect 22400 41331 22800 41337
rect 23400 41331 23800 41337
rect 2659 41277 4200 41282
rect 4600 41277 4829 41282
rect 21346 41326 23400 41331
rect 23800 41326 23922 41331
rect 4200 41271 4600 41277
rect 21346 41266 21351 41326
rect 21411 41266 21449 41326
rect 21509 41266 21749 41326
rect 21809 41266 22049 41326
rect 22109 41266 22349 41326
rect 22409 41266 22649 41326
rect 22709 41266 22949 41326
rect 23009 41266 23249 41326
rect 23309 41266 23400 41326
rect 23800 41266 23857 41326
rect 23917 41266 23922 41326
rect 21346 41261 23400 41266
rect 23800 41261 23922 41266
rect 21400 41255 21800 41261
rect 22400 41255 22800 41261
rect 23400 41255 23800 41261
rect 7800 40505 8200 40506
rect 8800 40505 9200 40506
rect 9800 40505 10200 40506
rect 13000 40505 13400 40506
rect 14000 40505 14400 40506
rect 15000 40505 15400 40506
rect 7739 40500 10327 40505
rect 7739 40430 7745 40500
rect 7815 40430 9800 40500
rect 10200 40430 10252 40500
rect 10322 40430 10327 40500
rect 7739 40425 10327 40430
rect 12939 40500 15527 40505
rect 12939 40430 12945 40500
rect 13015 40430 15000 40500
rect 15400 40430 15452 40500
rect 15522 40430 15527 40500
rect 12939 40425 15527 40430
rect 7800 40424 8200 40425
rect 8800 40424 9200 40425
rect 9800 40424 10200 40425
rect 13000 40424 13400 40425
rect 14000 40424 14400 40425
rect 15000 40424 15400 40425
rect 7800 40295 8200 40296
rect 8800 40295 9200 40296
rect 9800 40295 10200 40296
rect 13000 40295 13400 40296
rect 14000 40295 14400 40296
rect 15000 40295 15400 40296
rect 7711 40290 10347 40295
rect 7711 40220 7716 40290
rect 7786 40220 8800 40290
rect 9200 40220 10272 40290
rect 10342 40220 10347 40290
rect 3200 40215 3602 40220
rect 7711 40215 10347 40220
rect 12911 40290 15547 40295
rect 12911 40220 12916 40290
rect 12986 40220 14000 40290
rect 14400 40220 15472 40290
rect 15542 40220 15547 40290
rect 12911 40215 15547 40220
rect 2658 40214 4828 40215
rect 7800 40214 8200 40215
rect 8800 40214 9200 40215
rect 9800 40214 10200 40215
rect 13000 40214 13400 40215
rect 14000 40214 14400 40215
rect 15000 40214 15400 40215
rect 2658 40210 3200 40214
rect 3602 40210 4828 40214
rect 2658 40150 2663 40210
rect 2723 40150 2963 40210
rect 3023 40150 3200 40210
rect 3623 40150 3863 40210
rect 3923 40150 4163 40210
rect 4223 40150 4463 40210
rect 4523 40150 4763 40210
rect 4823 40150 4828 40210
rect 21400 40199 21800 40205
rect 22400 40199 22800 40205
rect 23400 40199 23800 40205
rect 2658 40145 3200 40150
rect 3602 40145 4828 40150
rect 21326 40194 22400 40199
rect 22800 40194 23952 40199
rect 3200 40138 3602 40144
rect 21326 40134 21331 40194
rect 21391 40134 21463 40194
rect 21523 40134 21763 40194
rect 21823 40134 22063 40194
rect 22123 40134 22363 40194
rect 22800 40134 22963 40194
rect 23023 40134 23263 40194
rect 23323 40134 23563 40194
rect 23623 40134 23887 40194
rect 23947 40134 23952 40194
rect 21326 40129 22400 40134
rect 22800 40129 23952 40134
rect 21400 40123 21800 40129
rect 22400 40123 22800 40129
rect 23400 40123 23800 40129
rect 7800 39163 8200 39164
rect 8800 39163 9200 39164
rect 9800 39163 10200 39164
rect 13000 39163 13400 39164
rect 14000 39163 14400 39164
rect 15000 39163 15400 39164
rect 7739 39158 10327 39163
rect 7739 39153 9800 39158
rect 10200 39153 10327 39158
rect 7739 39093 7751 39153
rect 7811 39093 8045 39153
rect 8105 39093 8345 39153
rect 8405 39093 8645 39153
rect 8705 39093 8945 39153
rect 9005 39093 9245 39153
rect 9305 39093 9545 39153
rect 9605 39093 9800 39153
rect 10205 39093 10257 39153
rect 10317 39093 10327 39153
rect 7739 39088 9800 39093
rect 10200 39088 10327 39093
rect 7739 39083 10327 39088
rect 12939 39158 15527 39163
rect 12939 39153 15000 39158
rect 15400 39153 15527 39158
rect 12939 39093 12951 39153
rect 13011 39093 13245 39153
rect 13305 39093 13545 39153
rect 13605 39093 13845 39153
rect 13905 39093 14145 39153
rect 14205 39093 14445 39153
rect 14505 39093 14745 39153
rect 14805 39093 15000 39153
rect 15405 39093 15457 39153
rect 15517 39093 15527 39153
rect 12939 39088 15000 39093
rect 15400 39088 15527 39093
rect 12939 39083 15527 39088
rect 7800 39082 8200 39083
rect 8800 39082 9200 39083
rect 9800 39082 10200 39083
rect 13000 39082 13400 39083
rect 14000 39082 14400 39083
rect 15000 39082 15400 39083
rect 21400 37838 21800 37844
rect 22400 37838 22800 37844
rect 23400 37838 23800 37844
rect 21346 37833 21400 37838
rect 21800 37833 23922 37838
rect 21346 37773 21351 37833
rect 21823 37773 22063 37833
rect 22123 37773 22363 37833
rect 22423 37773 22663 37833
rect 22723 37773 22963 37833
rect 23023 37773 23263 37833
rect 23323 37773 23563 37833
rect 23623 37773 23857 37833
rect 23917 37773 23922 37833
rect 21346 37768 21400 37773
rect 21800 37768 23922 37773
rect 21400 37762 21800 37768
rect 22400 37762 22800 37768
rect 23400 37762 23800 37768
rect 7800 36802 8200 36803
rect 8800 36802 9200 36803
rect 9800 36802 10200 36803
rect 13000 36802 13400 36803
rect 14000 36802 14400 36803
rect 15000 36802 15400 36803
rect 7711 36797 10347 36802
rect 7711 36792 8800 36797
rect 9200 36792 10347 36797
rect 7711 36732 7721 36792
rect 7781 36732 8045 36792
rect 8105 36732 8345 36792
rect 8405 36732 8645 36792
rect 8705 36732 8800 36792
rect 9200 36732 9245 36792
rect 9305 36732 9545 36792
rect 9605 36732 9845 36792
rect 9905 36732 10145 36792
rect 10205 36732 10277 36792
rect 10337 36732 10347 36792
rect 7711 36727 8800 36732
rect 9200 36727 10347 36732
rect 7711 36722 10347 36727
rect 12911 36797 15547 36802
rect 12911 36792 14000 36797
rect 14400 36792 15547 36797
rect 12911 36732 12921 36792
rect 12981 36732 13245 36792
rect 13305 36732 13545 36792
rect 13605 36732 13845 36792
rect 13905 36732 14000 36792
rect 14400 36732 14445 36792
rect 14505 36732 14745 36792
rect 14805 36732 15045 36792
rect 15105 36732 15345 36792
rect 15405 36732 15477 36792
rect 15537 36732 15547 36792
rect 12911 36727 14000 36732
rect 14400 36727 15547 36732
rect 12911 36722 15547 36727
rect 7800 36721 8200 36722
rect 8800 36721 9200 36722
rect 9800 36721 10200 36722
rect 13000 36721 13400 36722
rect 14000 36721 14400 36722
rect 15000 36721 15400 36722
rect 21400 36711 21800 36712
rect 22400 36711 22800 36712
rect 23400 36711 23800 36712
rect 21321 36706 23957 36711
rect 21321 36636 21326 36706
rect 21396 36636 22400 36706
rect 22800 36636 23882 36706
rect 23952 36636 23957 36706
rect 21321 36631 23957 36636
rect 21400 36630 21800 36631
rect 22400 36630 22800 36631
rect 23400 36630 23800 36631
rect 21400 36501 21800 36502
rect 22400 36501 22800 36502
rect 23400 36501 23800 36502
rect 21341 36496 23928 36501
rect 21341 36426 21346 36496
rect 21800 36426 23853 36496
rect 23923 36426 23928 36496
rect 21341 36421 23928 36426
rect 21400 36420 21800 36421
rect 22400 36420 22800 36421
rect 23400 36420 23800 36421
rect 7800 35670 8200 35671
rect 8800 35670 9200 35671
rect 9800 35670 10200 35671
rect 13000 35670 13400 35671
rect 14000 35670 14400 35671
rect 15000 35670 15400 35671
rect 7739 35665 10327 35670
rect 7739 35660 7800 35665
rect 8200 35660 10327 35665
rect 7739 35600 7751 35660
rect 8200 35600 8359 35660
rect 8419 35600 8659 35660
rect 8719 35600 8959 35660
rect 9019 35600 9259 35660
rect 9319 35600 9559 35660
rect 9619 35600 9859 35660
rect 9919 35600 10159 35660
rect 10219 35600 10257 35660
rect 10317 35600 10327 35660
rect 7739 35595 7800 35600
rect 8200 35595 10327 35600
rect 7739 35590 10327 35595
rect 12939 35665 15527 35670
rect 12939 35660 13000 35665
rect 13400 35660 15527 35665
rect 12939 35600 12951 35660
rect 13400 35600 13559 35660
rect 13619 35600 13859 35660
rect 13919 35600 14159 35660
rect 14219 35600 14459 35660
rect 14519 35600 14759 35660
rect 14819 35600 15059 35660
rect 15119 35600 15359 35660
rect 15419 35600 15457 35660
rect 15517 35600 15527 35660
rect 12939 35595 13000 35600
rect 13400 35595 15527 35600
rect 12939 35590 15527 35595
rect 7800 35589 8200 35590
rect 8800 35589 9200 35590
rect 9800 35589 10200 35590
rect 13000 35589 13400 35590
rect 14000 35589 14400 35590
rect 15000 35589 15400 35590
rect 21400 35369 21800 35370
rect 22400 35369 22800 35370
rect 23400 35369 23800 35370
rect 21321 35364 23957 35369
rect 21321 35359 22400 35364
rect 22800 35359 23957 35364
rect 21321 35299 21331 35359
rect 21391 35299 21462 35359
rect 21522 35299 21762 35359
rect 21822 35299 22062 35359
rect 22122 35299 22362 35359
rect 22800 35299 22962 35359
rect 23022 35299 23262 35359
rect 23322 35299 23562 35359
rect 23622 35299 23887 35359
rect 23947 35299 23957 35359
rect 21321 35294 22400 35299
rect 22800 35294 23957 35299
rect 21321 35289 23957 35294
rect 21400 35288 21800 35289
rect 22400 35288 22800 35289
rect 23400 35288 23800 35289
rect 7800 29209 8200 29215
rect 7784 29144 7800 29204
rect 8800 29204 9200 29215
rect 9800 29204 10200 29215
rect 13000 29209 13400 29215
rect 8200 29144 8217 29204
rect 8784 29144 9217 29204
rect 9784 29144 10217 29204
rect 12984 29144 13000 29204
rect 7800 29133 8200 29139
rect 8800 29133 9200 29144
rect 9800 29133 10200 29144
rect 14000 29204 14400 29215
rect 15000 29204 15400 29215
rect 13400 29144 13417 29204
rect 13984 29144 14417 29204
rect 14984 29144 15417 29204
rect 13000 29133 13400 29139
rect 14000 29133 14400 29144
rect 15000 29133 15400 29144
rect 7800 28833 8200 28915
rect 8800 28909 9200 28915
rect 8784 28844 8800 28904
rect 9800 28904 10200 28915
rect 13000 28904 13400 28915
rect 14000 28909 14400 28915
rect 9200 28844 9217 28904
rect 9784 28844 10217 28904
rect 12984 28844 13417 28904
rect 13984 28844 14000 28904
rect 8800 28833 9200 28839
rect 9800 28833 10200 28844
rect 13000 28833 13400 28844
rect 15000 28904 15400 28915
rect 14400 28844 14417 28904
rect 14984 28844 15417 28904
rect 14000 28833 14400 28839
rect 15000 28833 15400 28844
rect 7800 28609 8200 28615
rect 7784 28544 7800 28604
rect 8800 28604 9200 28615
rect 9800 28604 10200 28615
rect 13000 28609 13400 28615
rect 8200 28544 8217 28604
rect 8784 28544 9217 28604
rect 9784 28544 10217 28604
rect 12984 28544 13000 28604
rect 7800 28533 8200 28539
rect 8800 28533 9200 28544
rect 9800 28533 10200 28544
rect 14000 28604 14400 28615
rect 15000 28604 15400 28615
rect 13400 28544 13417 28604
rect 13984 28544 14417 28604
rect 14984 28544 15417 28604
rect 13000 28533 13400 28539
rect 14000 28533 14400 28544
rect 15000 28533 15400 28544
rect 7800 28304 8200 28315
rect 8800 28309 9200 28315
rect 7784 28244 8217 28304
rect 8784 28244 8800 28304
rect 7800 28233 8200 28244
rect 9800 28304 10200 28315
rect 13000 28304 13400 28315
rect 14000 28309 14400 28315
rect 9200 28244 9217 28304
rect 9784 28244 10217 28304
rect 12984 28244 13417 28304
rect 13984 28244 14000 28304
rect 8800 28233 9200 28239
rect 9800 28233 10200 28244
rect 13000 28233 13400 28244
rect 15000 28304 15400 28315
rect 14400 28244 14417 28304
rect 14984 28244 15417 28304
rect 14000 28233 14400 28239
rect 15000 28233 15400 28244
rect 7800 28009 8200 28015
rect 7784 27944 7800 28004
rect 8800 28004 9200 28015
rect 9800 28004 10200 28015
rect 13000 28009 13400 28015
rect 8200 27944 8217 28004
rect 8784 27944 9217 28004
rect 9784 27944 10217 28004
rect 12984 27944 13000 28004
rect 7800 27933 8200 27939
rect 8800 27933 9200 27944
rect 9800 27933 10200 27944
rect 14000 28004 14400 28015
rect 15000 28004 15400 28015
rect 13400 27944 13417 28004
rect 13984 27944 14417 28004
rect 14984 27944 15417 28004
rect 13000 27933 13400 27939
rect 14000 27933 14400 27944
rect 15000 27933 15400 27944
rect 7800 27704 8200 27715
rect 8800 27709 9200 27715
rect 7784 27644 8217 27704
rect 8784 27644 8800 27704
rect 7800 27633 8200 27644
rect 9800 27704 10200 27715
rect 13000 27704 13400 27715
rect 14000 27709 14400 27715
rect 9200 27644 9217 27704
rect 9784 27644 10217 27704
rect 12984 27644 13417 27704
rect 13984 27644 14000 27704
rect 8800 27633 9200 27639
rect 9800 27633 10200 27644
rect 13000 27633 13400 27644
rect 15000 27704 15400 27715
rect 14400 27644 14417 27704
rect 14984 27644 15417 27704
rect 14000 27633 14400 27639
rect 15000 27633 15400 27644
rect 7800 27409 8200 27415
rect 7784 27344 7800 27404
rect 8800 27404 9200 27415
rect 9800 27404 10200 27415
rect 13000 27409 13400 27415
rect 8200 27344 8217 27404
rect 8784 27344 9217 27404
rect 9784 27344 10217 27404
rect 12984 27344 13000 27404
rect 7800 27333 8200 27339
rect 8800 27333 9200 27344
rect 9800 27333 10200 27344
rect 14000 27404 14400 27415
rect 15000 27404 15400 27415
rect 13400 27344 13417 27404
rect 13984 27344 14417 27404
rect 14984 27344 15417 27404
rect 13000 27333 13400 27339
rect 14000 27333 14400 27344
rect 15000 27333 15400 27344
rect 7800 27104 8200 27115
rect 8800 27109 9200 27115
rect 7784 27044 8217 27104
rect 8784 27044 8800 27104
rect 7800 27033 8200 27044
rect 9800 27104 10200 27115
rect 13000 27104 13400 27115
rect 14000 27109 14400 27115
rect 9200 27044 9217 27104
rect 9784 27044 10217 27104
rect 12984 27044 13417 27104
rect 13984 27044 14000 27104
rect 8800 27033 9200 27039
rect 9800 27033 10200 27044
rect 13000 27033 13400 27044
rect 15000 27104 15400 27115
rect 14400 27044 14417 27104
rect 14984 27044 15417 27104
rect 14000 27033 14400 27039
rect 15000 27033 15400 27044
rect 7800 26809 8200 26815
rect 7784 26744 7800 26804
rect 8800 26804 9200 26815
rect 9800 26804 10200 26815
rect 13000 26809 13400 26815
rect 8200 26744 8217 26804
rect 8784 26744 9217 26804
rect 9784 26744 10217 26804
rect 12984 26744 13000 26804
rect 7800 26733 8200 26739
rect 8800 26733 9200 26744
rect 9800 26733 10200 26744
rect 14000 26804 14400 26815
rect 15000 26804 15400 26815
rect 13400 26744 13417 26804
rect 13984 26744 14417 26804
rect 14984 26744 15417 26804
rect 13000 26733 13400 26739
rect 14000 26733 14400 26744
rect 15000 26733 15400 26744
rect 21400 24600 21800 24606
rect 3200 24580 23800 24600
rect 3200 24220 7820 24580
rect 8180 24220 13020 24580
rect 13380 24220 21420 24580
rect 21780 24220 23800 24580
rect 3200 24200 23800 24220
rect 21400 24194 21800 24200
rect 3200 23600 3600 23606
rect 8800 23600 9200 23606
rect 3200 23580 23800 23600
rect 3200 23220 3220 23580
rect 3580 23220 8820 23580
rect 9180 23220 14020 23580
rect 14380 23220 22420 23580
rect 22780 23220 23800 23580
rect 3200 23200 23800 23220
rect 3200 23194 3600 23200
rect 8800 23194 9200 23200
rect 9800 22600 10200 22606
rect 15000 22600 15400 22606
rect 23400 22600 23800 22606
rect 3200 22580 23800 22600
rect 3200 22220 4220 22580
rect 4580 22220 9820 22580
rect 10180 22220 15020 22580
rect 15380 22220 23420 22580
rect 23780 22220 23800 22580
rect 3200 22200 23800 22220
rect 9800 22194 10200 22200
rect 15000 22194 15400 22200
rect 23400 22194 23800 22200
rect 7800 20602 8200 20608
rect 6895 20402 7800 20602
rect 8200 20402 9355 20602
rect 6895 6894 6955 20402
rect 7195 6654 7255 20162
rect 7495 6894 7555 20402
rect 7800 20396 8200 20402
rect 8095 20162 8155 20396
rect 7795 6654 7855 20162
rect 8087 6894 8093 20162
rect 8157 6894 8163 20162
rect 8395 6654 8455 20162
rect 8695 6894 8755 20402
rect 8987 6894 8993 20162
rect 9057 6894 9063 20162
rect 9295 6894 9355 20402
rect 13097 20008 13303 20014
rect 13097 19796 13303 19802
rect 14097 17422 14303 17428
rect 14097 17210 14303 17216
rect 13097 11003 13303 11009
rect 13097 10791 13303 10797
rect 14097 8015 14303 8021
rect 13688 7981 13836 7986
rect 13688 7843 13693 7981
rect 13831 7843 14097 7981
rect 13688 7838 13836 7843
rect 14097 7803 14303 7809
rect 8997 6660 9057 6894
rect 13000 6719 13400 6725
rect 21400 6719 21800 6725
rect 8800 6654 9200 6660
rect 7195 6454 8800 6654
rect 13400 6519 21400 6719
rect 13000 6513 13400 6519
rect 8800 6448 9200 6454
rect 17323 6419 17523 6519
rect 21400 6513 21800 6519
rect 17323 6281 17354 6419
rect 17492 6281 17523 6419
rect 17323 6250 17523 6281
rect 14000 5069 14400 5075
rect 22400 5069 22800 5075
rect 13522 4869 14000 5069
rect 14400 4869 22400 5069
rect 14000 4863 14400 4869
rect 17323 4595 17523 4869
rect 22400 4863 22797 4869
rect 17323 4457 17354 4595
rect 17492 4457 17523 4595
rect 17323 4426 17523 4457
<< via3 >>
rect 8800 41627 9200 41632
rect 8800 41567 8946 41627
rect 8946 41567 9006 41627
rect 9006 41567 9200 41627
rect 8800 41562 9200 41567
rect 14000 41627 14400 41632
rect 14000 41567 14146 41627
rect 14146 41567 14206 41627
rect 14206 41567 14400 41627
rect 14000 41562 14400 41567
rect 4200 41342 4600 41347
rect 4200 41282 4224 41342
rect 4224 41282 4464 41342
rect 4464 41282 4524 41342
rect 4524 41282 4600 41342
rect 4200 41277 4600 41282
rect 23400 41326 23800 41331
rect 23400 41266 23549 41326
rect 23549 41266 23609 41326
rect 23609 41266 23800 41326
rect 23400 41261 23800 41266
rect 9800 40430 10200 40500
rect 15000 40430 15400 40500
rect 8800 40220 9200 40290
rect 14000 40220 14400 40290
rect 3200 40210 3602 40214
rect 3200 40150 3263 40210
rect 3263 40150 3323 40210
rect 3323 40150 3563 40210
rect 3563 40150 3602 40210
rect 3200 40144 3602 40150
rect 22400 40194 22800 40199
rect 22400 40134 22423 40194
rect 22423 40134 22663 40194
rect 22663 40134 22723 40194
rect 22723 40134 22800 40194
rect 22400 40129 22800 40134
rect 9800 39153 10200 39158
rect 9800 39093 9845 39153
rect 9845 39093 9905 39153
rect 9905 39093 10145 39153
rect 10145 39093 10200 39153
rect 9800 39088 10200 39093
rect 15000 39153 15400 39158
rect 15000 39093 15045 39153
rect 15045 39093 15105 39153
rect 15105 39093 15345 39153
rect 15345 39093 15400 39153
rect 15000 39088 15400 39093
rect 21400 37833 21800 37838
rect 21400 37773 21411 37833
rect 21411 37773 21463 37833
rect 21463 37773 21523 37833
rect 21523 37773 21763 37833
rect 21763 37773 21800 37833
rect 21400 37768 21800 37773
rect 8800 36792 9200 36797
rect 8800 36732 8945 36792
rect 8945 36732 9005 36792
rect 9005 36732 9200 36792
rect 8800 36727 9200 36732
rect 14000 36792 14400 36797
rect 14000 36732 14145 36792
rect 14145 36732 14205 36792
rect 14205 36732 14400 36792
rect 14000 36727 14400 36732
rect 22400 36636 22800 36706
rect 21400 36426 21416 36496
rect 21416 36426 21800 36496
rect 7800 35660 8200 35665
rect 7800 35600 7811 35660
rect 7811 35600 8059 35660
rect 8059 35600 8119 35660
rect 8119 35600 8200 35660
rect 7800 35595 8200 35600
rect 13000 35660 13400 35665
rect 13000 35600 13011 35660
rect 13011 35600 13259 35660
rect 13259 35600 13319 35660
rect 13319 35600 13400 35660
rect 13000 35595 13400 35600
rect 22400 35359 22800 35364
rect 22400 35299 22422 35359
rect 22422 35299 22662 35359
rect 22662 35299 22722 35359
rect 22722 35299 22800 35359
rect 22400 35294 22800 35299
rect 7800 29139 8200 29209
rect 13000 29139 13400 29209
rect 8800 28839 9200 28909
rect 14000 28839 14400 28909
rect 7800 28539 8200 28609
rect 13000 28539 13400 28609
rect 8800 28239 9200 28309
rect 14000 28239 14400 28309
rect 7800 27939 8200 28009
rect 13000 27939 13400 28009
rect 8800 27639 9200 27709
rect 14000 27639 14400 27709
rect 7800 27339 8200 27409
rect 13000 27339 13400 27409
rect 8800 27039 9200 27109
rect 14000 27039 14400 27109
rect 7800 26739 8200 26809
rect 13000 26739 13400 26809
rect 7820 24220 8180 24580
rect 13020 24220 13380 24580
rect 21420 24220 21780 24580
rect 3220 23220 3580 23580
rect 8820 23220 9180 23580
rect 14020 23220 14380 23580
rect 22420 23220 22780 23580
rect 4220 22220 4580 22580
rect 9820 22220 10180 22580
rect 15020 22220 15380 22580
rect 23420 22220 23780 22580
rect 7800 20402 8200 20602
rect 8093 6894 8157 20162
rect 8993 6894 9057 20162
rect 13097 19974 13303 20008
rect 13097 19836 13131 19974
rect 13131 19836 13269 19974
rect 13269 19836 13303 19974
rect 13097 19802 13303 19836
rect 14097 17388 14303 17422
rect 14097 17250 14131 17388
rect 14131 17250 14269 17388
rect 14269 17250 14303 17388
rect 14097 17216 14303 17250
rect 13097 10969 13303 11003
rect 13097 10831 13131 10969
rect 13131 10831 13269 10969
rect 13269 10831 13303 10969
rect 13097 10797 13303 10831
rect 14097 7809 14303 8015
rect 8800 6454 9200 6654
rect 13000 6519 13400 6719
rect 21400 6519 21800 6719
rect 14000 4869 14400 5069
rect 22400 4869 22800 5069
<< metal4 >>
rect 3200 40215 3600 44152
rect 4200 41348 4600 44152
rect 7800 41633 8200 44152
rect 8800 41633 9200 44152
rect 9800 41633 10200 44152
rect 13000 41633 13400 44152
rect 14000 41633 14400 44152
rect 15000 41633 15400 44152
rect 7799 41561 8201 41633
rect 8799 41632 9201 41633
rect 8799 41562 8800 41632
rect 9200 41562 9201 41632
rect 8799 41561 9201 41562
rect 9799 41561 10201 41633
rect 12999 41561 13401 41633
rect 13999 41632 14401 41633
rect 13999 41562 14000 41632
rect 14400 41562 14401 41632
rect 13999 41561 14401 41562
rect 14999 41561 15401 41633
rect 4199 41347 4601 41348
rect 4199 41277 4200 41347
rect 4600 41277 4601 41347
rect 4199 41276 4601 41277
rect 3199 40214 3603 40215
rect 3199 40144 3200 40214
rect 3602 40144 3603 40214
rect 3199 40143 3603 40144
rect 3200 23601 3600 40143
rect 3199 23580 3601 23601
rect 3199 23220 3220 23580
rect 3580 23220 3601 23580
rect 3199 23199 3601 23220
rect 3200 1000 3600 23199
rect 4200 22601 4600 41276
rect 7800 40501 8200 41561
rect 8800 40501 9200 41561
rect 9800 40501 10200 41561
rect 13000 40501 13400 41561
rect 14000 40501 14400 41561
rect 15000 40501 15400 41561
rect 21400 41332 21800 44152
rect 22400 41332 22800 44152
rect 23400 41332 23800 44152
rect 21399 41260 21801 41332
rect 22399 41260 22801 41332
rect 23399 41331 23801 41332
rect 23399 41261 23400 41331
rect 23800 41261 23801 41331
rect 23399 41260 23801 41261
rect 7799 40429 8201 40501
rect 8799 40429 9201 40501
rect 9799 40500 10201 40501
rect 9799 40430 9800 40500
rect 10200 40430 10201 40500
rect 9799 40429 10201 40430
rect 12999 40429 13401 40501
rect 13999 40429 14401 40501
rect 14999 40500 15401 40501
rect 14999 40430 15000 40500
rect 15400 40430 15401 40500
rect 14999 40429 15401 40430
rect 7800 40291 8200 40429
rect 8800 40291 9200 40429
rect 9800 40291 10200 40429
rect 13000 40291 13400 40429
rect 14000 40291 14400 40429
rect 15000 40291 15400 40429
rect 7799 40219 8201 40291
rect 8799 40290 9201 40291
rect 8799 40220 8800 40290
rect 9200 40220 9201 40290
rect 8799 40219 9201 40220
rect 9799 40219 10201 40291
rect 12999 40219 13401 40291
rect 13999 40290 14401 40291
rect 13999 40220 14000 40290
rect 14400 40220 14401 40290
rect 13999 40219 14401 40220
rect 14999 40219 15401 40291
rect 7800 39159 8200 40219
rect 8800 39159 9200 40219
rect 9800 39159 10200 40219
rect 13000 39159 13400 40219
rect 14000 39159 14400 40219
rect 15000 39159 15400 40219
rect 21400 40200 21800 41260
rect 22400 40200 22800 41260
rect 23400 40200 23800 41260
rect 21399 40128 21801 40200
rect 22399 40199 22801 40200
rect 22399 40129 22400 40199
rect 22800 40129 22801 40199
rect 22399 40128 22801 40129
rect 23399 40128 23801 40200
rect 7799 39087 8201 39159
rect 8799 39087 9201 39159
rect 9799 39158 10201 39159
rect 9799 39088 9800 39158
rect 10200 39088 10201 39158
rect 9799 39087 10201 39088
rect 12999 39087 13401 39159
rect 13999 39087 14401 39159
rect 14999 39158 15401 39159
rect 14999 39088 15000 39158
rect 15400 39088 15401 39158
rect 14999 39087 15401 39088
rect 7800 36798 8200 39087
rect 8800 36798 9200 39087
rect 9800 36798 10200 39087
rect 13000 36798 13400 39087
rect 14000 36798 14400 39087
rect 15000 36798 15400 39087
rect 21400 37839 21800 40128
rect 22400 37839 22800 40128
rect 23400 37839 23800 40128
rect 21399 37838 21801 37839
rect 21399 37768 21400 37838
rect 21800 37768 21801 37838
rect 21399 37767 21801 37768
rect 22399 37767 22801 37839
rect 23399 37767 23801 37839
rect 7799 36726 8201 36798
rect 8799 36797 9201 36798
rect 8799 36727 8800 36797
rect 9200 36727 9201 36797
rect 8799 36726 9201 36727
rect 9799 36726 10201 36798
rect 12999 36726 13401 36798
rect 13999 36797 14401 36798
rect 13999 36727 14000 36797
rect 14400 36727 14401 36797
rect 13999 36726 14401 36727
rect 14999 36726 15401 36798
rect 7800 35666 8200 36726
rect 8800 35666 9200 36726
rect 9800 35666 10200 36726
rect 13000 35666 13400 36726
rect 14000 35666 14400 36726
rect 15000 35666 15400 36726
rect 21400 36707 21800 37767
rect 22400 36707 22800 37767
rect 23400 36707 23800 37767
rect 21399 36635 21801 36707
rect 22399 36706 22801 36707
rect 22399 36636 22400 36706
rect 22800 36636 22801 36706
rect 22399 36635 22801 36636
rect 23399 36635 23801 36707
rect 21400 36497 21800 36635
rect 22400 36497 22800 36635
rect 23400 36497 23800 36635
rect 21399 36496 21801 36497
rect 21399 36426 21400 36496
rect 21800 36426 21801 36496
rect 21399 36425 21801 36426
rect 22399 36425 22801 36497
rect 23399 36425 23801 36497
rect 7799 35665 8201 35666
rect 7799 35595 7800 35665
rect 8200 35595 8201 35665
rect 7799 35594 8201 35595
rect 8799 35594 9201 35666
rect 9799 35594 10201 35666
rect 12999 35665 13401 35666
rect 12999 35595 13000 35665
rect 13400 35595 13401 35665
rect 12999 35594 13401 35595
rect 13999 35594 14401 35666
rect 14999 35594 15401 35666
rect 7800 35456 8200 35594
rect 8800 35456 9200 35594
rect 9800 35456 10200 35594
rect 7799 35384 8201 35456
rect 8799 35384 9201 35456
rect 9799 35384 10201 35456
rect 7800 29210 8200 35384
rect 8800 29210 9200 35384
rect 9800 29210 10200 35384
rect 13000 29210 13400 35594
rect 14000 29210 14400 35594
rect 15000 29210 15400 35594
rect 21400 35365 21800 36425
rect 22400 35365 22800 36425
rect 23400 35365 23800 36425
rect 21399 35293 21801 35365
rect 22399 35364 22801 35365
rect 22399 35294 22400 35364
rect 22800 35294 22801 35364
rect 22399 35293 22801 35294
rect 23399 35293 23801 35365
rect 7799 29209 8201 29210
rect 7799 29139 7800 29209
rect 8200 29139 8201 29209
rect 7799 29138 8201 29139
rect 8799 29138 9201 29210
rect 9799 29138 10201 29210
rect 12999 29209 13401 29210
rect 12999 29139 13000 29209
rect 13400 29139 13401 29209
rect 12999 29138 13401 29139
rect 13999 29138 14401 29210
rect 14999 29138 15401 29210
rect 7800 28910 8200 29138
rect 8800 28910 9200 29138
rect 9800 28910 10200 29138
rect 13000 28910 13400 29138
rect 14000 28910 14400 29138
rect 15000 28910 15400 29138
rect 7799 28838 8201 28910
rect 8799 28909 9201 28910
rect 8799 28839 8800 28909
rect 9200 28839 9201 28909
rect 8799 28838 9201 28839
rect 9799 28838 10201 28910
rect 12999 28838 13401 28910
rect 13999 28909 14401 28910
rect 13999 28839 14000 28909
rect 14400 28839 14401 28909
rect 13999 28838 14401 28839
rect 14999 28838 15401 28910
rect 7800 28610 8200 28838
rect 8800 28610 9200 28838
rect 9800 28610 10200 28838
rect 13000 28610 13400 28838
rect 14000 28610 14400 28838
rect 15000 28610 15400 28838
rect 7799 28609 8201 28610
rect 7799 28539 7800 28609
rect 8200 28539 8201 28609
rect 7799 28538 8201 28539
rect 8799 28538 9201 28610
rect 9799 28538 10201 28610
rect 12999 28609 13401 28610
rect 12999 28539 13000 28609
rect 13400 28539 13401 28609
rect 12999 28538 13401 28539
rect 13999 28538 14401 28610
rect 14999 28538 15401 28610
rect 7800 28310 8200 28538
rect 8800 28310 9200 28538
rect 9800 28310 10200 28538
rect 13000 28310 13400 28538
rect 14000 28310 14400 28538
rect 15000 28310 15400 28538
rect 7799 28238 8201 28310
rect 8799 28309 9201 28310
rect 8799 28239 8800 28309
rect 9200 28239 9201 28309
rect 8799 28238 9201 28239
rect 9799 28238 10201 28310
rect 12999 28238 13401 28310
rect 13999 28309 14401 28310
rect 13999 28239 14000 28309
rect 14400 28239 14401 28309
rect 13999 28238 14401 28239
rect 14999 28238 15401 28310
rect 7800 28010 8200 28238
rect 8800 28010 9200 28238
rect 9800 28010 10200 28238
rect 13000 28010 13400 28238
rect 14000 28010 14400 28238
rect 15000 28010 15400 28238
rect 7799 28009 8201 28010
rect 7799 27939 7800 28009
rect 8200 27939 8201 28009
rect 7799 27938 8201 27939
rect 8799 27938 9201 28010
rect 9799 27938 10201 28010
rect 12999 28009 13401 28010
rect 12999 27939 13000 28009
rect 13400 27939 13401 28009
rect 12999 27938 13401 27939
rect 13999 27938 14401 28010
rect 14999 27938 15401 28010
rect 7800 27710 8200 27938
rect 8800 27710 9200 27938
rect 9800 27710 10200 27938
rect 13000 27710 13400 27938
rect 14000 27710 14400 27938
rect 15000 27710 15400 27938
rect 7799 27638 8201 27710
rect 8799 27709 9201 27710
rect 8799 27639 8800 27709
rect 9200 27639 9201 27709
rect 8799 27638 9201 27639
rect 9799 27638 10201 27710
rect 12999 27638 13401 27710
rect 13999 27709 14401 27710
rect 13999 27639 14000 27709
rect 14400 27639 14401 27709
rect 13999 27638 14401 27639
rect 14999 27638 15401 27710
rect 7800 27410 8200 27638
rect 8800 27410 9200 27638
rect 9800 27410 10200 27638
rect 13000 27410 13400 27638
rect 14000 27410 14400 27638
rect 15000 27410 15400 27638
rect 7799 27409 8201 27410
rect 7799 27339 7800 27409
rect 8200 27339 8201 27409
rect 7799 27338 8201 27339
rect 8799 27338 9201 27410
rect 9799 27338 10201 27410
rect 12999 27409 13401 27410
rect 12999 27339 13000 27409
rect 13400 27339 13401 27409
rect 12999 27338 13401 27339
rect 13999 27338 14401 27410
rect 14999 27338 15401 27410
rect 7800 27110 8200 27338
rect 8800 27110 9200 27338
rect 9800 27110 10200 27338
rect 13000 27110 13400 27338
rect 14000 27110 14400 27338
rect 15000 27110 15400 27338
rect 7799 27038 8201 27110
rect 8799 27109 9201 27110
rect 8799 27039 8800 27109
rect 9200 27039 9201 27109
rect 8799 27038 9201 27039
rect 9799 27038 10201 27110
rect 12999 27038 13401 27110
rect 13999 27109 14401 27110
rect 13999 27039 14000 27109
rect 14400 27039 14401 27109
rect 13999 27038 14401 27039
rect 14999 27038 15401 27110
rect 7800 26810 8200 27038
rect 8800 26810 9200 27038
rect 9800 26810 10200 27038
rect 13000 26810 13400 27038
rect 14000 26810 14400 27038
rect 15000 26810 15400 27038
rect 7799 26809 8201 26810
rect 7799 26739 7800 26809
rect 8200 26739 8201 26809
rect 7799 26738 8201 26739
rect 8799 26738 9201 26810
rect 9799 26738 10201 26810
rect 12999 26809 13401 26810
rect 12999 26739 13000 26809
rect 13400 26739 13401 26809
rect 12999 26738 13401 26739
rect 13999 26738 14401 26810
rect 14999 26738 15401 26810
rect 7800 24601 8200 26738
rect 7799 24580 8201 24601
rect 7799 24220 7820 24580
rect 8180 24220 8201 24580
rect 7799 24199 8201 24220
rect 4199 22580 4601 22601
rect 4199 22220 4220 22580
rect 4580 22220 4601 22580
rect 4199 22199 4601 22220
rect 4200 1000 4600 22199
rect 7800 20603 8200 24199
rect 8800 23601 9200 26738
rect 8799 23580 9201 23601
rect 8799 23220 8820 23580
rect 9180 23220 9201 23580
rect 8799 23199 9201 23220
rect 7799 20602 8201 20603
rect 7799 20402 7800 20602
rect 8200 20402 8201 20602
rect 7799 20401 8201 20402
rect 7800 20162 8200 20401
rect 7800 6894 8093 20162
rect 8157 6894 8200 20162
rect 7800 1000 8200 6894
rect 8800 20162 9200 23199
rect 9800 22601 10200 26738
rect 13000 24601 13400 26738
rect 12999 24580 13401 24601
rect 12999 24220 13020 24580
rect 13380 24220 13401 24580
rect 12999 24199 13401 24220
rect 9799 22580 10201 22601
rect 9799 22220 9820 22580
rect 10180 22220 10201 22580
rect 9799 22199 10201 22220
rect 8800 6894 8993 20162
rect 9057 6894 9200 20162
rect 8800 6655 9200 6894
rect 8799 6654 9201 6655
rect 8799 6454 8800 6654
rect 9200 6454 9201 6654
rect 8799 6453 9201 6454
rect 8800 1000 9200 6453
rect 9800 1000 10200 22199
rect 13000 20008 13400 24199
rect 14000 23601 14400 26738
rect 13999 23580 14401 23601
rect 13999 23220 14020 23580
rect 14380 23220 14401 23580
rect 13999 23199 14401 23220
rect 13000 19802 13097 20008
rect 13303 19802 13400 20008
rect 13000 11003 13400 19802
rect 13000 10797 13097 11003
rect 13303 10797 13400 11003
rect 13000 6720 13400 10797
rect 14000 17457 14400 23199
rect 15000 22601 15400 26738
rect 21400 24601 21800 35293
rect 21399 24580 21801 24601
rect 21399 24220 21420 24580
rect 21780 24220 21801 24580
rect 21399 24199 21801 24220
rect 14999 22580 15401 22601
rect 14999 22220 15020 22580
rect 15380 22220 15401 22580
rect 14999 22199 15401 22220
rect 14000 17422 14401 17457
rect 14000 17216 14097 17422
rect 14303 17216 14401 17422
rect 14000 17181 14401 17216
rect 14000 8015 14400 17181
rect 14000 7809 14097 8015
rect 14303 7809 14400 8015
rect 12999 6719 13401 6720
rect 12999 6519 13000 6719
rect 13400 6519 13401 6719
rect 12999 6518 13401 6519
rect 13000 1000 13400 6518
rect 14000 5070 14400 7809
rect 13999 5069 14401 5070
rect 13999 4869 14000 5069
rect 14400 4869 14401 5069
rect 13999 4868 14401 4869
rect 14000 1000 14400 4868
rect 15000 1000 15400 22199
rect 21400 6720 21800 24199
rect 22400 23601 22800 35293
rect 22399 23580 22801 23601
rect 22399 23220 22420 23580
rect 22780 23220 22801 23580
rect 22399 23199 22801 23220
rect 21399 6719 21801 6720
rect 21399 6519 21400 6719
rect 21800 6519 21801 6719
rect 21399 6518 21801 6519
rect 21400 1000 21800 6518
rect 22400 5070 22800 23199
rect 23400 22601 23800 35293
rect 23399 22580 23801 22601
rect 23399 22220 23420 22580
rect 23780 22220 23801 22580
rect 23399 22199 23801 22220
rect 22399 5069 22801 5070
rect 22399 4869 22400 5069
rect 22800 4869 22801 5069
rect 22399 4868 22801 4869
rect 22400 1000 22800 4868
rect 23400 1000 23800 22199
<< labels >>
flabel metal4 7800 1000 8200 44152 1 FreeSans 400 0 0 0 VAPWR
port 0 nsew power bidirectional
flabel metal4 8800 1000 9200 44152 1 FreeSans 400 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 9800 1000 10200 44152 1 FreeSans 400 0 0 0 VDPWR
port 1 nsew power bidirectional
flabel metal4 13000 1000 13400 44152 1 FreeSans 400 0 0 0 VAPWR
port 0 nsew power bidirectional
flabel metal4 14000 1000 14400 44152 1 FreeSans 400 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 15000 1000 15400 44152 1 FreeSans 400 0 0 0 VDPWR
port 1 nsew power bidirectional
flabel metal4 21400 1000 21800 44152 1 FreeSans 400 0 0 0 VAPWR
port 0 nsew power bidirectional
flabel metal4 22400 1000 22800 44152 1 FreeSans 400 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 23400 1000 23800 44152 1 FreeSans 400 0 0 0 VDPWR
port 1 nsew power bidirectional
flabel metal4 3200 1000 3600 44152 1 FreeSans 400 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 4200 1000 4600 44152 1 FreeSans 400 0 0 0 VDPWR
port 1 nsew power bidirectional
<< end >>
