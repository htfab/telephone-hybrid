magic
tech sky130A
magscale 1 2
timestamp 1731100676
<< metal1 >>
rect 276 3473 346 3490
rect 276 3076 285 3473
rect 337 3076 346 3473
rect 276 3058 346 3076
rect 1438 3058 1674 3490
rect 3578 2648 3716 2654
rect 3578 2504 3716 2510
rect 3854 1436 3992 1442
rect 3854 1292 3992 1298
rect 2340 767 2532 773
rect 2340 715 2352 767
rect 2520 715 2532 767
rect 2340 709 2532 715
rect 2716 767 2908 773
rect 2716 715 2728 767
rect 2896 715 2908 767
rect 2716 709 2908 715
<< via1 >>
rect 285 3076 337 3473
rect 3578 2510 3716 2648
rect 3854 1298 3992 1436
rect 2352 715 2520 767
rect 2728 715 2896 767
<< metal2 >>
rect 277 12216 415 12354
rect 6990 4605 7867 4639
rect 276 3473 346 3490
rect 276 3106 285 3473
rect 121 3076 285 3106
rect 337 3076 346 3473
rect 6990 3263 7867 3297
rect 121 3058 346 3076
rect 121 917 169 3058
rect 3392 2714 3483 2762
rect 3290 2236 3350 2245
rect 3290 2167 3350 2176
rect 276 985 414 1123
rect 3296 917 3344 2167
rect 121 869 2460 917
rect 2412 773 2460 869
rect 2788 869 3344 917
rect 2788 773 2836 869
rect 3392 821 3440 2714
rect 3572 2510 3578 2648
rect 3716 2510 3722 2648
rect 3076 773 3440 821
rect 2340 767 2532 773
rect 2340 715 2352 767
rect 2520 715 2532 767
rect 2340 709 2532 715
rect 2716 767 2908 773
rect 2716 715 2728 767
rect 2896 715 2908 767
rect 2716 709 2908 715
rect 3076 -1033 3124 773
rect 3578 -175 3716 2510
rect 6990 1921 7867 1955
rect 3848 1298 3854 1436
rect 3992 1298 3998 1436
rect 3574 -303 3583 -175
rect 3711 -303 3720 -175
rect 3578 -308 3716 -303
rect 2914 -1081 3124 -1033
rect 110 -1733 310 -1533
rect 3854 -1825 3992 1298
rect 6990 579 7867 613
rect 3850 -1953 3859 -1825
rect 3987 -1953 3996 -1825
rect 110 -2249 310 -2049
<< via2 >>
rect 3290 2176 3350 2236
rect 3583 -303 3711 -175
rect 3859 -1953 3987 -1825
<< metal3 >>
rect 3285 2236 3355 2241
rect 2625 2176 3290 2236
rect 3350 2176 3355 2236
rect 3285 2171 3355 2176
rect 2811 -175 3716 -170
rect 2811 -303 3583 -175
rect 3711 -303 3716 -175
rect 2811 -308 3716 -303
rect 2811 -1825 3992 -1820
rect 2811 -1953 3859 -1825
rect 3987 -1953 3992 -1825
rect 2811 -1958 3992 -1953
use opamp  x1
timestamp 1727597281
transform 1 0 -3094 0 1 -827
box 3204 -1676 6132 1720
use digipot  x2
timestamp 1731100676
transform 1 0 0 0 1 943
box 110 -943 7867 12467
<< labels >>
flabel metal1 1438 3058 1674 3490 0 FreeSans 128 0 0 0 IN
port 4 nsew
flabel metal2 110 -2249 310 -2049 0 FreeSans 128 0 0 0 OUT
port 6 nsew
flabel metal2 110 -1733 310 -1533 0 FreeSans 128 0 0 0 LINE
port 5 nsew
flabel metal2 277 12216 415 12354 0 FreeSans 128 0 0 0 VDD
port 7 nsew
flabel metal2 276 985 414 1123 0 FreeSans 128 0 0 0 VSS
port 8 nsew
flabel metal2 6990 579 7867 613 0 FreeSans 128 0 0 0 D3
port 3 nsew
flabel metal2 6990 1921 7867 1955 0 FreeSans 128 0 0 0 D0
port 0 nsew
flabel metal2 6990 3263 7867 3297 0 FreeSans 128 0 0 0 D1
port 1 nsew
flabel metal2 6990 4605 7867 4639 0 FreeSans 128 0 0 0 D2
port 2 nsew
<< end >>
