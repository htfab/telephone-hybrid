magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< dnwell >>
rect -365 -275 4076 10803
<< nwell >>
rect -445 10597 4156 10883
rect -445 -69 -159 10597
rect 3870 -69 4156 10597
rect -445 -355 4156 -69
<< nsubdiff >>
rect -408 10826 4119 10846
rect -408 10792 -328 10826
rect 4039 10792 4119 10826
rect -408 10772 4119 10792
rect -408 10766 -334 10772
rect -408 -238 -388 10766
rect -354 -238 -334 10766
rect -408 -244 -334 -238
rect 4045 10766 4119 10772
rect 4045 -238 4065 10766
rect 4099 -238 4119 10766
rect 4045 -244 4119 -238
rect -408 -264 4119 -244
rect -408 -298 -328 -264
rect 4039 -298 4119 -264
rect -408 -318 4119 -298
<< nsubdiffcont >>
rect -328 10792 4039 10826
rect -388 -238 -354 10766
rect 4065 -238 4099 10766
rect -328 -298 4039 -264
<< locali >>
rect -388 10792 -328 10826
rect 4039 10792 4099 10826
rect -388 10766 -354 10792
rect -388 -264 -354 -238
rect 4065 10766 4099 10792
rect 4065 -264 4099 -238
rect -388 -298 -328 -264
rect 4039 -298 4099 -264
use hybrid  hybrid_0
timestamp 1727597281
transform 1 0 -3204 0 1 3276
box 3204 -3276 7092 7391
<< end >>
