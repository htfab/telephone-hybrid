magic
tech sky130A
magscale 1 2
timestamp 1727641872
<< metal1 >>
rect 0 44952 200 45152
rect 28872 44952 29072 45152
rect 0 0 200 200
rect 28872 0 29072 200
use decoder4_signed_dnwell  decoder4_signed_dnwell_0
timestamp 1727641872
transform 0 -1 18656 1 0 26230
box -381 -415 3987 14056
use hybrid_ctrl_dnwell  hybrid_ctrl_dnwell_0
timestamp 1727641872
transform -1 0 13998 0 1 4355
box -686 -355 7998 16559
use hybrid_dnwell  hybrid_dnwell_0
timestamp 1727597281
transform 1 0 20445 0 1 4355
box -445 -355 4156 10883
use passgate_dnwell  passgate_dnwell_0
timestamp 1727641355
transform 1 0 17134 0 1 4415
box -734 -415 1210 2762
use shifters_dnwell  shifters_dnwell_0
timestamp 1727641773
transform -1 0 10382 0 -1 41662
box -686 -415 3382 6813
use shifters_dnwell  shifters_dnwell_2
timestamp 1727641773
transform -1 0 15582 0 -1 41662
box -686 -415 3382 6813
use shifters_dnwell  shifters_dnwell_3
timestamp 1727641773
transform 1 0 21286 0 1 35264
box -686 -415 3382 6813
use signal_routing  signal_routing_0
timestamp 1727631305
transform 1 0 0 0 1 0
box 0 0 29072 45152
use tie_highs_dnwell  tie_highs_dnwell_0
timestamp 1727641773
transform 1 0 2486 0 1 40115
box -686 -415 3382 1978
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
