magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< error_p >>
rect -144 166 144 200
rect -186 -166 186 166
rect -144 -200 144 -166
<< nwell >>
rect -144 -200 144 200
<< mvpmos >>
rect -50 -100 50 100
<< mvpdiff >>
rect -120 88 -50 100
rect -120 -88 -108 88
rect -74 -88 -50 88
rect -120 -100 -50 -88
rect 50 88 120 100
rect 50 -88 74 88
rect 108 -88 120 88
rect 50 -100 120 -88
<< mvpdiffc >>
rect -108 -88 -74 88
rect 74 -88 108 88
<< poly >>
rect -50 181 50 197
rect -50 147 -34 181
rect 34 147 50 181
rect -50 100 50 147
rect -50 -147 50 -100
rect -50 -181 -34 -147
rect 34 -181 50 -147
rect -50 -197 50 -181
<< polycont >>
rect -34 147 34 181
rect -34 -181 34 -147
<< locali >>
rect -50 147 -34 181
rect 34 147 50 181
rect -108 88 -74 104
rect -108 -104 -74 -88
rect 74 88 108 104
rect 74 -104 108 -88
rect -50 -181 -34 -147
rect 34 -181 50 -147
<< viali >>
rect -34 147 34 181
rect -108 -88 -74 88
rect 74 -88 108 88
rect -34 -181 34 -147
<< metal1 >>
rect -46 181 46 187
rect -46 147 -34 181
rect 34 147 46 181
rect -46 141 46 147
rect -114 88 -68 100
rect -114 -88 -108 88
rect -74 -88 -68 88
rect -114 -100 -68 -88
rect 68 88 114 100
rect 68 -88 74 88
rect 108 -88 114 88
rect 68 -100 114 -88
rect -46 -147 46 -141
rect -46 -181 -34 -147
rect 34 -181 46 -147
rect -46 -187 46 -181
<< end >>
