magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< error_p >>
rect -108 109 -50 239
rect 50 109 108 239
rect -108 -239 -50 -109
rect 50 -239 108 -109
<< mvnmos >>
rect -50 109 50 239
rect -50 -239 50 -109
<< mvndiff >>
rect -108 227 -50 239
rect -108 121 -96 227
rect -62 121 -50 227
rect -108 109 -50 121
rect 50 227 108 239
rect 50 121 62 227
rect 96 121 108 227
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -227 -96 -121
rect -62 -227 -50 -121
rect -108 -239 -50 -227
rect 50 -121 108 -109
rect 50 -227 62 -121
rect 96 -227 108 -121
rect 50 -239 108 -227
<< mvndiffc >>
rect -96 121 -62 227
rect 62 121 96 227
rect -96 -227 -62 -121
rect 62 -227 96 -121
<< poly >>
rect -50 311 50 327
rect -50 277 -34 311
rect 34 277 50 311
rect -50 239 50 277
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -277 50 -239
rect -50 -311 -34 -277
rect 34 -311 50 -277
rect -50 -327 50 -311
<< polycont >>
rect -34 277 34 311
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -311 34 -277
<< locali >>
rect -50 277 -34 311
rect 34 277 50 311
rect -96 227 -62 243
rect -96 105 -62 121
rect 62 227 96 243
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -243 -62 -227
rect 62 -121 96 -105
rect 62 -243 96 -227
rect -50 -311 -34 -277
rect 34 -311 50 -277
<< viali >>
rect -34 277 34 311
rect -96 121 -62 227
rect 62 121 96 227
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -227 -62 -121
rect 62 -227 96 -121
rect -34 -311 34 -277
<< metal1 >>
rect -46 311 46 317
rect -46 277 -34 311
rect 34 277 46 311
rect -46 271 46 277
rect -102 227 -56 239
rect -102 121 -96 227
rect -62 121 -56 227
rect -102 109 -56 121
rect 56 227 102 239
rect 56 121 62 227
rect 96 121 102 227
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -227 -96 -121
rect -62 -227 -56 -121
rect -102 -239 -56 -227
rect 56 -121 102 -109
rect 56 -227 62 -121
rect 96 -227 102 -121
rect 56 -239 102 -227
rect -46 -277 46 -271
rect -46 -311 -34 -277
rect 34 -311 46 -277
rect -46 -317 46 -311
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.65 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
