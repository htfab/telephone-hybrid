magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< xpolycontact >>
rect -616 3184 -546 3616
rect -616 -3616 -546 -3184
rect -450 3184 -380 3616
rect -450 -3616 -380 -3184
rect -284 3184 -214 3616
rect -284 -3616 -214 -3184
rect -118 3184 -48 3616
rect -118 -3616 -48 -3184
rect 48 3184 118 3616
rect 48 -3616 118 -3184
rect 214 3184 284 3616
rect 214 -3616 284 -3184
rect 380 3184 450 3616
rect 380 -3616 450 -3184
rect 546 3184 616 3616
rect 546 -3616 616 -3184
<< xpolyres >>
rect -616 -3184 -546 3184
rect -450 -3184 -380 3184
rect -284 -3184 -214 3184
rect -118 -3184 -48 3184
rect 48 -3184 118 3184
rect 214 -3184 284 3184
rect 380 -3184 450 3184
rect 546 -3184 616 3184
<< viali >>
rect -600 3201 -562 3598
rect -434 3201 -396 3598
rect -268 3201 -230 3598
rect -102 3201 -64 3598
rect 64 3201 102 3598
rect 230 3201 268 3598
rect 396 3201 434 3598
rect 562 3201 600 3598
rect -600 -3598 -562 -3201
rect -434 -3598 -396 -3201
rect -268 -3598 -230 -3201
rect -102 -3598 -64 -3201
rect 64 -3598 102 -3201
rect 230 -3598 268 -3201
rect 396 -3598 434 -3201
rect 562 -3598 600 -3201
<< metal1 >>
rect -606 3598 -556 3610
rect -606 3201 -600 3598
rect -562 3201 -556 3598
rect -606 3189 -556 3201
rect -440 3598 -390 3610
rect -440 3201 -434 3598
rect -396 3201 -390 3598
rect -440 3189 -390 3201
rect -274 3598 -224 3610
rect -274 3201 -268 3598
rect -230 3201 -224 3598
rect -274 3189 -224 3201
rect -108 3598 -58 3610
rect -108 3201 -102 3598
rect -64 3201 -58 3598
rect -108 3189 -58 3201
rect 58 3598 108 3610
rect 58 3201 64 3598
rect 102 3201 108 3598
rect 58 3189 108 3201
rect 224 3598 274 3610
rect 224 3201 230 3598
rect 268 3201 274 3598
rect 224 3189 274 3201
rect 390 3598 440 3610
rect 390 3201 396 3598
rect 434 3201 440 3598
rect 390 3189 440 3201
rect 556 3598 606 3610
rect 556 3201 562 3598
rect 600 3201 606 3598
rect 556 3189 606 3201
rect -606 -3201 -556 -3189
rect -606 -3598 -600 -3201
rect -562 -3598 -556 -3201
rect -606 -3610 -556 -3598
rect -440 -3201 -390 -3189
rect -440 -3598 -434 -3201
rect -396 -3598 -390 -3201
rect -440 -3610 -390 -3598
rect -274 -3201 -224 -3189
rect -274 -3598 -268 -3201
rect -230 -3598 -224 -3201
rect -274 -3610 -224 -3598
rect -108 -3201 -58 -3189
rect -108 -3598 -102 -3201
rect -64 -3598 -58 -3201
rect -108 -3610 -58 -3598
rect 58 -3201 108 -3189
rect 58 -3598 64 -3201
rect 102 -3598 108 -3201
rect 58 -3610 108 -3598
rect 224 -3201 274 -3189
rect 224 -3598 230 -3201
rect 268 -3598 274 -3201
rect 224 -3610 274 -3598
rect 390 -3201 440 -3189
rect 390 -3598 396 -3201
rect 434 -3598 440 -3201
rect 390 -3610 440 -3598
rect 556 -3201 606 -3189
rect 556 -3598 562 -3201
rect 600 -3598 606 -3201
rect 556 -3610 606 -3598
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 32 m 1 nx 8 wmin 0.350 lmin 0.50 rho 2000 val 183.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
