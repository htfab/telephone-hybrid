magic
tech sky130A
timestamp 1727597281
<< nwell >>
rect -30 303 94 646
<< pwell >>
rect -25 0 94 278
<< mvpsubdiff >>
rect -7 231 44 260
rect -7 206 22 231
rect -7 72 -1 206
rect 16 72 22 206
rect -7 47 22 72
rect -7 18 44 47
<< mvnsubdiff >>
rect 3 584 44 613
rect 3 559 32 584
rect 3 390 9 559
rect 26 390 32 559
rect 3 365 32 390
rect 3 336 44 365
<< mvpsubdiffcont >>
rect -1 72 16 206
<< mvnsubdiffcont >>
rect 9 390 26 559
<< locali >>
rect 9 590 44 607
rect 9 559 26 590
rect 9 359 26 390
rect 9 342 44 359
rect -1 237 44 254
rect -1 206 16 237
rect -1 41 16 72
rect -1 24 44 41
<< end >>
