magic
tech sky130A
magscale 1 2
timestamp 1731100676
<< dnwell >>
rect -606 -275 8058 16479
<< nwell >>
rect -686 16273 8138 16559
rect -686 -69 -400 16273
rect 7852 -69 8138 16273
rect -686 -355 8138 -69
<< nsubdiff >>
rect -649 16502 8101 16522
rect -649 16468 -569 16502
rect 8021 16468 8101 16502
rect -649 16448 8101 16468
rect -649 16442 -575 16448
rect -649 -238 -629 16442
rect -595 -238 -575 16442
rect -649 -244 -575 -238
rect 8027 16442 8101 16448
rect 8027 -238 8047 16442
rect 8081 -238 8101 16442
rect 8027 -244 8101 -238
rect -649 -264 8101 -244
rect -649 -298 -569 -264
rect 8021 -298 8101 -264
rect -649 -318 8101 -298
<< nsubdiffcont >>
rect -569 16468 8021 16502
rect -629 -238 -595 16442
rect 8047 -238 8081 16442
rect -569 -298 8021 -264
<< locali >>
rect -629 16468 -569 16502
rect 8021 16468 8081 16502
rect -629 16442 -595 16468
rect -629 -264 -595 -238
rect 8047 16442 8081 16468
rect 8047 -264 8081 -238
rect -629 -298 -569 -264
rect 8021 -298 8081 -264
use hybrid_ctrl  hybrid_ctrl_0
timestamp 1731100676
transform 1 0 -110 0 1 2503
box 110 -2503 7867 13410
<< end >>
