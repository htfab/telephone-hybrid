magic
tech sky130A
magscale 1 2
timestamp 1727641872
<< dnwell >>
rect -606 -275 7918 16479
<< nwell >>
rect -686 16273 7998 16559
rect -686 -69 -400 16273
rect 7712 -69 7998 16273
rect -686 -355 7998 -69
<< nsubdiff >>
rect -649 16502 7961 16522
rect -649 16468 -569 16502
rect 7881 16468 7961 16502
rect -649 16448 7961 16468
rect -649 16442 -575 16448
rect -649 -238 -629 16442
rect -595 -238 -575 16442
rect -649 -244 -575 -238
rect 7887 16442 7961 16448
rect 7887 -238 7907 16442
rect 7941 -238 7961 16442
rect 7887 -244 7961 -238
rect -649 -264 7961 -244
rect -649 -298 -569 -264
rect 7881 -298 7961 -264
rect -649 -318 7961 -298
<< nsubdiffcont >>
rect -569 16468 7881 16502
rect -629 -238 -595 16442
rect 7907 -238 7941 16442
rect -569 -298 7881 -264
<< locali >>
rect -629 16468 -569 16502
rect 7881 16468 7941 16502
rect -629 16442 -595 16468
rect -629 -264 -595 -238
rect 7907 16442 7941 16468
rect 7907 -264 7941 -238
rect -629 -298 -569 -264
rect 7881 -298 7941 -264
use hybrid_ctrl  hybrid_ctrl_0
timestamp 1727641872
transform 1 0 -110 0 1 2503
box 110 -2503 7727 13410
<< end >>
