magic
tech sky130A
magscale 1 2
timestamp 1727641178
<< metal2 >>
rect 166 1866 2788 2004
rect 268 1193 406 1601
rect 2752 1193 2890 1601
rect 166 180 304 685
rect 452 557 570 675
rect 728 557 846 675
rect 1004 557 1122 675
rect 1280 557 1398 675
rect 1556 557 1674 675
rect 1832 557 1950 675
rect 2108 557 2226 675
rect 2384 557 2502 675
rect 2650 180 2788 685
rect 166 42 2788 180
<< via2 >>
rect 554 1203 672 1321
rect 830 1203 948 1321
rect 1106 1203 1224 1321
rect 1382 1203 1500 1321
rect 1658 1203 1776 1321
rect 1934 1203 2052 1321
rect 2210 1203 2328 1321
rect 2486 1203 2604 1321
<< metal3 >>
rect 544 1321 2614 1331
rect 544 1203 554 1321
rect 672 1203 830 1321
rect 948 1203 1106 1321
rect 1224 1203 1382 1321
rect 1500 1203 1658 1321
rect 1776 1203 1934 1321
rect 2052 1203 2210 1321
rect 2328 1203 2486 1321
rect 2604 1203 2614 1321
rect 544 1193 2614 1203
rect 622 1192 682 1193
rect 898 1192 958 1193
rect 1174 1192 1234 1193
rect 1450 1192 1510 1193
rect 1726 1192 1786 1193
rect 2002 1192 2062 1193
rect 2278 1192 2338 1193
rect 2554 1192 2614 1193
use transistor_quartet_bus10  transistor_quartet_bus10_0
timestamp 1727641178
transform 1 0 0 0 1 0
box 0 0 3056 2076
use passgate  x1
timestamp 1727641004
transform 1 0 324 0 1 0
box 112 42 358 2004
use passgate  x2
timestamp 1727641004
transform 1 0 600 0 1 0
box 112 42 358 2004
use passgate  x3
timestamp 1727641004
transform 1 0 876 0 1 0
box 112 42 358 2004
use passgate  x4
timestamp 1727641004
transform 1 0 1152 0 1 0
box 112 42 358 2004
use passgate  x5
timestamp 1727641004
transform 1 0 1428 0 1 0
box 112 42 358 2004
use passgate  x6
timestamp 1727641004
transform 1 0 1704 0 1 0
box 112 42 358 2004
use passgate  x7
timestamp 1727641004
transform 1 0 1980 0 1 0
box 112 42 358 2004
use passgate  x8
timestamp 1727641004
transform 1 0 2256 0 1 0
box 112 42 358 2004
use passgate  xdummy1
timestamp 1727641004
transform 1 0 48 0 1 0
box 112 42 358 2004
use passgate  xdummy2
timestamp 1727641004
transform 1 0 2532 0 1 0
box 112 42 358 2004
<< end >>
