magic
tech sky130A
magscale 1 2
timestamp 1727637843
<< nwell >>
rect -60 606 2636 1292
<< pwell >>
rect -60 556 126 557
rect -60 0 2636 556
<< mvnmos >>
rect 188 213 288 343
rect 488 213 588 343
rect 788 213 888 343
rect 1088 213 1188 343
rect 1388 213 1488 343
rect 1688 213 1788 343
rect 1988 213 2088 343
rect 2288 213 2388 343
<< mvpmos >>
rect 188 849 288 1049
rect 488 849 588 1049
rect 788 849 888 1049
rect 1088 849 1188 1049
rect 1388 849 1488 1049
rect 1688 849 1788 1049
rect 1988 849 2088 1049
rect 2288 849 2388 1049
<< mvndiff >>
rect 118 331 188 343
rect 118 225 130 331
rect 164 225 188 331
rect 118 213 188 225
rect 288 331 358 343
rect 288 225 312 331
rect 346 225 358 331
rect 288 213 358 225
rect 418 331 488 343
rect 418 225 430 331
rect 464 225 488 331
rect 418 213 488 225
rect 588 331 658 343
rect 588 225 612 331
rect 646 225 658 331
rect 588 213 658 225
rect 718 331 788 343
rect 718 225 730 331
rect 764 225 788 331
rect 718 213 788 225
rect 888 331 958 343
rect 888 225 912 331
rect 946 225 958 331
rect 888 213 958 225
rect 1018 331 1088 343
rect 1018 225 1030 331
rect 1064 225 1088 331
rect 1018 213 1088 225
rect 1188 331 1258 343
rect 1188 225 1212 331
rect 1246 225 1258 331
rect 1188 213 1258 225
rect 1318 331 1388 343
rect 1318 225 1330 331
rect 1364 225 1388 331
rect 1318 213 1388 225
rect 1488 331 1558 343
rect 1488 225 1512 331
rect 1546 225 1558 331
rect 1488 213 1558 225
rect 1618 331 1688 343
rect 1618 225 1630 331
rect 1664 225 1688 331
rect 1618 213 1688 225
rect 1788 331 1858 343
rect 1788 225 1812 331
rect 1846 225 1858 331
rect 1788 213 1858 225
rect 1918 331 1988 343
rect 1918 225 1930 331
rect 1964 225 1988 331
rect 1918 213 1988 225
rect 2088 331 2158 343
rect 2088 225 2112 331
rect 2146 225 2158 331
rect 2088 213 2158 225
rect 2218 331 2288 343
rect 2218 225 2230 331
rect 2264 225 2288 331
rect 2218 213 2288 225
rect 2388 331 2458 343
rect 2388 225 2412 331
rect 2446 225 2458 331
rect 2388 213 2458 225
<< mvpdiff >>
rect 118 1037 188 1049
rect 118 861 130 1037
rect 164 861 188 1037
rect 118 849 188 861
rect 288 1037 358 1049
rect 288 861 312 1037
rect 346 861 358 1037
rect 288 849 358 861
rect 418 1037 488 1049
rect 418 861 430 1037
rect 464 861 488 1037
rect 418 849 488 861
rect 588 1037 658 1049
rect 588 861 612 1037
rect 646 861 658 1037
rect 588 849 658 861
rect 718 1037 788 1049
rect 718 861 730 1037
rect 764 861 788 1037
rect 718 849 788 861
rect 888 1037 958 1049
rect 888 861 912 1037
rect 946 861 958 1037
rect 888 849 958 861
rect 1018 1037 1088 1049
rect 1018 861 1030 1037
rect 1064 861 1088 1037
rect 1018 849 1088 861
rect 1188 1037 1258 1049
rect 1188 861 1212 1037
rect 1246 861 1258 1037
rect 1188 849 1258 861
rect 1318 1037 1388 1049
rect 1318 861 1330 1037
rect 1364 861 1388 1037
rect 1318 849 1388 861
rect 1488 1037 1558 1049
rect 1488 861 1512 1037
rect 1546 861 1558 1037
rect 1488 849 1558 861
rect 1618 1037 1688 1049
rect 1618 861 1630 1037
rect 1664 861 1688 1037
rect 1618 849 1688 861
rect 1788 1037 1858 1049
rect 1788 861 1812 1037
rect 1846 861 1858 1037
rect 1788 849 1858 861
rect 1918 1037 1988 1049
rect 1918 861 1930 1037
rect 1964 861 1988 1037
rect 1918 849 1988 861
rect 2088 1037 2158 1049
rect 2088 861 2112 1037
rect 2146 861 2158 1037
rect 2088 849 2158 861
rect 2218 1037 2288 1049
rect 2218 861 2230 1037
rect 2264 861 2288 1037
rect 2218 849 2288 861
rect 2388 1037 2458 1049
rect 2388 861 2412 1037
rect 2446 861 2458 1037
rect 2388 849 2458 861
<< mvndiffc >>
rect 130 225 164 331
rect 312 225 346 331
rect 430 225 464 331
rect 612 225 646 331
rect 730 225 764 331
rect 912 225 946 331
rect 1030 225 1064 331
rect 1212 225 1246 331
rect 1330 225 1364 331
rect 1512 225 1546 331
rect 1630 225 1664 331
rect 1812 225 1846 331
rect 1930 225 1964 331
rect 2112 225 2146 331
rect 2230 225 2264 331
rect 2412 225 2446 331
<< mvpdiffc >>
rect 130 861 164 1037
rect 312 861 346 1037
rect 430 861 464 1037
rect 612 861 646 1037
rect 730 861 764 1037
rect 912 861 946 1037
rect 1030 861 1064 1037
rect 1212 861 1246 1037
rect 1330 861 1364 1037
rect 1512 861 1546 1037
rect 1630 861 1664 1037
rect 1812 861 1846 1037
rect 1930 861 1964 1037
rect 2112 861 2146 1037
rect 2230 861 2264 1037
rect 2412 861 2446 1037
<< mvpsubdiff >>
rect -14 508 2600 520
rect -14 474 124 508
rect 352 474 424 508
rect 652 474 724 508
rect 952 474 1024 508
rect 1252 474 1324 508
rect 1552 474 1624 508
rect 1852 474 1924 508
rect 2152 474 2224 508
rect 2452 474 2600 508
rect -14 462 2600 474
rect -14 412 44 462
rect -14 144 -2 412
rect 32 144 44 412
rect 2542 412 2600 462
rect -14 94 44 144
rect 2542 144 2554 412
rect 2588 144 2600 412
rect 2542 94 2600 144
rect -14 82 2600 94
rect -14 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2600 82
rect -14 36 2600 48
<< mvnsubdiff >>
rect 6 1214 2570 1226
rect 6 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2570 1214
rect 6 1168 2570 1180
rect 6 1118 64 1168
rect 6 780 18 1118
rect 52 780 64 1118
rect 2512 1118 2570 1168
rect 6 730 64 780
rect 2512 780 2524 1118
rect 2558 780 2570 1118
rect 2512 730 2570 780
rect 6 718 2570 730
rect 6 684 124 718
rect 352 684 424 718
rect 652 684 724 718
rect 952 684 1024 718
rect 1252 684 1324 718
rect 1552 684 1624 718
rect 1852 684 1924 718
rect 2152 684 2224 718
rect 2452 684 2570 718
rect 6 672 2570 684
<< mvpsubdiffcont >>
rect 124 474 352 508
rect 424 474 652 508
rect 724 474 952 508
rect 1024 474 1252 508
rect 1324 474 1552 508
rect 1624 474 1852 508
rect 1924 474 2152 508
rect 2224 474 2452 508
rect -2 144 32 412
rect 2554 144 2588 412
rect 124 48 352 82
rect 424 48 652 82
rect 724 48 952 82
rect 1024 48 1252 82
rect 1324 48 1552 82
rect 1624 48 1852 82
rect 1924 48 2152 82
rect 2224 48 2452 82
<< mvnsubdiffcont >>
rect 124 1180 352 1214
rect 424 1180 652 1214
rect 724 1180 952 1214
rect 1024 1180 1252 1214
rect 1324 1180 1552 1214
rect 1624 1180 1852 1214
rect 1924 1180 2152 1214
rect 2224 1180 2452 1214
rect 18 780 52 1118
rect 2524 780 2558 1118
rect 124 684 352 718
rect 424 684 652 718
rect 724 684 952 718
rect 1024 684 1252 718
rect 1324 684 1552 718
rect 1624 684 1852 718
rect 1924 684 2152 718
rect 2224 684 2452 718
<< poly >>
rect 188 1130 288 1146
rect 188 1096 204 1130
rect 272 1096 288 1130
rect 188 1049 288 1096
rect 488 1130 588 1146
rect 488 1096 504 1130
rect 572 1096 588 1130
rect 488 1049 588 1096
rect 788 1130 888 1146
rect 788 1096 804 1130
rect 872 1096 888 1130
rect 788 1049 888 1096
rect 1088 1130 1188 1146
rect 1088 1096 1104 1130
rect 1172 1096 1188 1130
rect 1088 1049 1188 1096
rect 1388 1130 1488 1146
rect 1388 1096 1404 1130
rect 1472 1096 1488 1130
rect 1388 1049 1488 1096
rect 1688 1130 1788 1146
rect 1688 1096 1704 1130
rect 1772 1096 1788 1130
rect 1688 1049 1788 1096
rect 1988 1130 2088 1146
rect 1988 1096 2004 1130
rect 2072 1096 2088 1130
rect 1988 1049 2088 1096
rect 2288 1130 2388 1146
rect 2288 1096 2304 1130
rect 2372 1096 2388 1130
rect 2288 1049 2388 1096
rect 188 802 288 849
rect 188 768 204 802
rect 272 768 288 802
rect 188 752 288 768
rect 488 802 588 849
rect 488 768 504 802
rect 572 768 588 802
rect 488 752 588 768
rect 788 802 888 849
rect 788 768 804 802
rect 872 768 888 802
rect 788 752 888 768
rect 1088 802 1188 849
rect 1088 768 1104 802
rect 1172 768 1188 802
rect 1088 752 1188 768
rect 1388 802 1488 849
rect 1388 768 1404 802
rect 1472 768 1488 802
rect 1388 752 1488 768
rect 1688 802 1788 849
rect 1688 768 1704 802
rect 1772 768 1788 802
rect 1688 752 1788 768
rect 1988 802 2088 849
rect 1988 768 2004 802
rect 2072 768 2088 802
rect 1988 752 2088 768
rect 2288 802 2388 849
rect 2288 768 2304 802
rect 2372 768 2388 802
rect 2288 752 2388 768
rect 188 415 288 431
rect 188 381 204 415
rect 272 381 288 415
rect 188 343 288 381
rect 488 415 588 431
rect 488 381 504 415
rect 572 381 588 415
rect 488 343 588 381
rect 788 415 888 431
rect 788 381 804 415
rect 872 381 888 415
rect 788 343 888 381
rect 1088 415 1188 431
rect 1088 381 1104 415
rect 1172 381 1188 415
rect 1088 343 1188 381
rect 1388 415 1488 431
rect 1388 381 1404 415
rect 1472 381 1488 415
rect 1388 343 1488 381
rect 1688 415 1788 431
rect 1688 381 1704 415
rect 1772 381 1788 415
rect 1688 343 1788 381
rect 1988 415 2088 431
rect 1988 381 2004 415
rect 2072 381 2088 415
rect 1988 343 2088 381
rect 2288 415 2388 431
rect 2288 381 2304 415
rect 2372 381 2388 415
rect 2288 343 2388 381
rect 188 175 288 213
rect 188 141 204 175
rect 272 141 288 175
rect 188 125 288 141
rect 488 175 588 213
rect 488 141 504 175
rect 572 141 588 175
rect 488 125 588 141
rect 788 175 888 213
rect 788 141 804 175
rect 872 141 888 175
rect 788 125 888 141
rect 1088 175 1188 213
rect 1088 141 1104 175
rect 1172 141 1188 175
rect 1088 125 1188 141
rect 1388 175 1488 213
rect 1388 141 1404 175
rect 1472 141 1488 175
rect 1388 125 1488 141
rect 1688 175 1788 213
rect 1688 141 1704 175
rect 1772 141 1788 175
rect 1688 125 1788 141
rect 1988 175 2088 213
rect 1988 141 2004 175
rect 2072 141 2088 175
rect 1988 125 2088 141
rect 2288 175 2388 213
rect 2288 141 2304 175
rect 2372 141 2388 175
rect 2288 125 2388 141
<< polycont >>
rect 204 1096 272 1130
rect 504 1096 572 1130
rect 804 1096 872 1130
rect 1104 1096 1172 1130
rect 1404 1096 1472 1130
rect 1704 1096 1772 1130
rect 2004 1096 2072 1130
rect 2304 1096 2372 1130
rect 204 768 272 802
rect 504 768 572 802
rect 804 768 872 802
rect 1104 768 1172 802
rect 1404 768 1472 802
rect 1704 768 1772 802
rect 2004 768 2072 802
rect 2304 768 2372 802
rect 204 381 272 415
rect 504 381 572 415
rect 804 381 872 415
rect 1104 381 1172 415
rect 1404 381 1472 415
rect 1704 381 1772 415
rect 2004 381 2072 415
rect 2304 381 2372 415
rect 204 141 272 175
rect 504 141 572 175
rect 804 141 872 175
rect 1104 141 1172 175
rect 1404 141 1472 175
rect 1704 141 1772 175
rect 2004 141 2072 175
rect 2304 141 2372 175
<< locali >>
rect 18 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2558 1214
rect 18 1118 52 1180
rect 188 1096 204 1130
rect 272 1096 288 1130
rect 488 1096 504 1130
rect 572 1096 588 1130
rect 788 1096 804 1130
rect 872 1096 888 1130
rect 1088 1096 1104 1130
rect 1172 1096 1188 1130
rect 1388 1096 1404 1130
rect 1472 1096 1488 1130
rect 1688 1096 1704 1130
rect 1772 1096 1788 1130
rect 1988 1096 2004 1130
rect 2072 1096 2088 1130
rect 2288 1096 2304 1130
rect 2372 1096 2388 1130
rect 2524 1118 2558 1180
rect 130 1037 164 1053
rect 130 845 164 861
rect 312 1037 346 1053
rect 312 845 346 861
rect 430 1037 464 1053
rect 430 845 464 861
rect 612 1037 646 1053
rect 612 845 646 861
rect 730 1037 764 1053
rect 730 845 764 861
rect 912 1037 946 1053
rect 912 845 946 861
rect 1030 1037 1064 1053
rect 1030 845 1064 861
rect 1212 1037 1246 1053
rect 1212 845 1246 861
rect 1330 1037 1364 1053
rect 1330 845 1364 861
rect 1512 1037 1546 1053
rect 1512 845 1546 861
rect 1630 1037 1664 1053
rect 1630 845 1664 861
rect 1812 1037 1846 1053
rect 1812 845 1846 861
rect 1930 1037 1964 1053
rect 1930 845 1964 861
rect 2112 1037 2146 1053
rect 2112 845 2146 861
rect 2230 1037 2264 1053
rect 2230 845 2264 861
rect 2412 1037 2446 1053
rect 2412 845 2446 861
rect 18 718 52 780
rect 188 768 204 802
rect 272 768 288 802
rect 488 768 504 802
rect 572 768 588 802
rect 788 768 804 802
rect 872 768 888 802
rect 1088 768 1104 802
rect 1172 768 1188 802
rect 1388 768 1404 802
rect 1472 768 1488 802
rect 1688 768 1704 802
rect 1772 768 1788 802
rect 1988 768 2004 802
rect 2072 768 2088 802
rect 2288 768 2304 802
rect 2372 768 2388 802
rect 2524 718 2558 780
rect 18 684 124 718
rect 352 684 424 718
rect 652 684 724 718
rect 952 684 1024 718
rect 1252 684 1324 718
rect 1552 684 1624 718
rect 1852 684 1924 718
rect 2152 684 2224 718
rect 2452 684 2558 718
rect -2 474 124 508
rect 352 474 424 508
rect 652 474 724 508
rect 952 474 1024 508
rect 1252 474 1324 508
rect 1552 474 1624 508
rect 1852 474 1924 508
rect 2152 474 2224 508
rect 2452 474 2588 508
rect -2 412 32 474
rect 188 381 204 415
rect 272 381 288 415
rect 488 381 504 415
rect 572 381 588 415
rect 788 381 804 415
rect 872 381 888 415
rect 1088 381 1104 415
rect 1172 381 1188 415
rect 1388 381 1404 415
rect 1472 381 1488 415
rect 1688 381 1704 415
rect 1772 381 1788 415
rect 1988 381 2004 415
rect 2072 381 2088 415
rect 2288 381 2304 415
rect 2372 381 2388 415
rect 2554 412 2588 474
rect 130 331 164 347
rect 130 209 164 225
rect 312 331 346 347
rect 312 209 346 225
rect 430 331 464 347
rect 430 209 464 225
rect 612 331 646 347
rect 612 209 646 225
rect 730 331 764 347
rect 730 209 764 225
rect 912 331 946 347
rect 912 209 946 225
rect 1030 331 1064 347
rect 1030 209 1064 225
rect 1212 331 1246 347
rect 1212 209 1246 225
rect 1330 331 1364 347
rect 1330 209 1364 225
rect 1512 331 1546 347
rect 1512 209 1546 225
rect 1630 331 1664 347
rect 1630 209 1664 225
rect 1812 331 1846 347
rect 1812 209 1846 225
rect 1930 331 1964 347
rect 1930 209 1964 225
rect 2112 331 2146 347
rect 2112 209 2146 225
rect 2230 331 2264 347
rect 2230 209 2264 225
rect 2412 331 2446 347
rect 2412 209 2446 225
rect -2 82 32 144
rect 188 141 204 175
rect 272 141 288 175
rect 488 141 504 175
rect 572 141 588 175
rect 788 141 804 175
rect 872 141 888 175
rect 1088 141 1104 175
rect 1172 141 1188 175
rect 1388 141 1404 175
rect 1472 141 1488 175
rect 1688 141 1704 175
rect 1772 141 1788 175
rect 1988 141 2004 175
rect 2072 141 2088 175
rect 2288 141 2304 175
rect 2372 141 2388 175
rect 2554 82 2588 144
rect -2 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2588 82
<< viali >>
rect 124 1180 352 1214
rect 424 1180 652 1214
rect 724 1180 952 1214
rect 1024 1180 1252 1214
rect 1324 1180 1552 1214
rect 1624 1180 1852 1214
rect 1924 1180 2152 1214
rect 2224 1180 2452 1214
rect 204 1096 272 1130
rect 504 1096 572 1130
rect 804 1096 872 1130
rect 1104 1096 1172 1130
rect 1404 1096 1472 1130
rect 1704 1096 1772 1130
rect 2004 1096 2072 1130
rect 2304 1096 2372 1130
rect 130 861 164 1037
rect 312 861 346 1037
rect 430 861 464 1037
rect 612 861 646 1037
rect 730 861 764 1037
rect 912 861 946 1037
rect 1030 861 1064 1037
rect 1212 861 1246 1037
rect 1330 861 1364 1037
rect 1512 861 1546 1037
rect 1630 861 1664 1037
rect 1812 861 1846 1037
rect 1930 861 1964 1037
rect 2112 861 2146 1037
rect 2230 861 2264 1037
rect 2412 861 2446 1037
rect 204 768 272 802
rect 504 768 572 802
rect 804 768 872 802
rect 1104 768 1172 802
rect 1404 768 1472 802
rect 1704 768 1772 802
rect 2004 768 2072 802
rect 2304 768 2372 802
rect 204 381 272 415
rect 504 381 572 415
rect 804 381 872 415
rect 1104 381 1172 415
rect 1404 381 1472 415
rect 1704 381 1772 415
rect 2004 381 2072 415
rect 2304 381 2372 415
rect 130 225 164 331
rect 312 225 346 331
rect 430 225 464 331
rect 612 225 646 331
rect 730 225 764 331
rect 912 225 946 331
rect 1030 225 1064 331
rect 1212 225 1246 331
rect 1330 225 1364 331
rect 1512 225 1546 331
rect 1630 225 1664 331
rect 1812 225 1846 331
rect 1930 225 1964 331
rect 2112 225 2146 331
rect 2230 225 2264 331
rect 2412 225 2446 331
rect 204 141 272 175
rect 504 141 572 175
rect 804 141 872 175
rect 1104 141 1172 175
rect 1404 141 1472 175
rect 1704 141 1772 175
rect 2004 141 2072 175
rect 2304 141 2372 175
rect 124 48 352 82
rect 424 48 652 82
rect 724 48 952 82
rect 1024 48 1252 82
rect 1324 48 1552 82
rect 1624 48 1852 82
rect 1924 48 2152 82
rect 2224 48 2452 82
<< metal1 >>
rect 88 1214 2488 1226
rect 88 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2488 1214
rect 88 1168 2488 1180
rect 192 1130 284 1136
rect 192 1096 204 1130
rect 272 1096 284 1130
rect 192 1090 284 1096
rect 492 1130 584 1136
rect 492 1096 504 1130
rect 572 1096 584 1130
rect 492 1090 584 1096
rect 792 1130 884 1136
rect 792 1096 804 1130
rect 872 1096 884 1130
rect 792 1090 884 1096
rect 1092 1130 1184 1136
rect 1092 1096 1104 1130
rect 1172 1096 1184 1130
rect 1092 1090 1184 1096
rect 1392 1130 1484 1136
rect 1392 1096 1404 1130
rect 1472 1096 1484 1130
rect 1392 1090 1484 1096
rect 1692 1130 1784 1136
rect 1692 1096 1704 1130
rect 1772 1096 1784 1130
rect 1692 1090 1784 1096
rect 1992 1130 2084 1136
rect 1992 1096 2004 1130
rect 2072 1096 2084 1130
rect 1992 1090 2084 1096
rect 2292 1130 2384 1136
rect 2292 1096 2304 1130
rect 2372 1096 2384 1130
rect 2292 1090 2384 1096
rect 130 1049 164 1053
rect 124 1037 170 1049
rect 124 861 130 1037
rect 164 861 170 1037
rect 124 849 170 861
rect 130 845 164 849
rect 221 808 255 1090
rect 312 1049 346 1053
rect 430 1049 464 1053
rect 306 1037 352 1049
rect 306 861 312 1037
rect 346 861 352 1037
rect 306 849 352 861
rect 424 1037 470 1049
rect 424 861 430 1037
rect 464 861 470 1037
rect 424 849 470 861
rect 312 845 346 849
rect 430 845 464 849
rect 521 808 555 1090
rect 612 1049 646 1053
rect 730 1049 764 1053
rect 606 1037 652 1049
rect 606 861 612 1037
rect 646 861 652 1037
rect 606 849 652 861
rect 724 1037 770 1049
rect 724 861 730 1037
rect 764 861 770 1037
rect 724 849 770 861
rect 612 845 646 849
rect 730 845 764 849
rect 821 808 855 1090
rect 912 1049 946 1053
rect 1030 1049 1064 1053
rect 906 1037 952 1049
rect 906 861 912 1037
rect 946 861 952 1037
rect 906 849 952 861
rect 1024 1037 1070 1049
rect 1024 861 1030 1037
rect 1064 861 1070 1037
rect 1024 849 1070 861
rect 912 845 946 849
rect 1030 845 1064 849
rect 1121 808 1155 1090
rect 1212 1049 1246 1053
rect 1330 1049 1364 1053
rect 1206 1037 1252 1049
rect 1206 861 1212 1037
rect 1246 861 1252 1037
rect 1206 849 1252 861
rect 1324 1037 1370 1049
rect 1324 861 1330 1037
rect 1364 861 1370 1037
rect 1324 849 1370 861
rect 1212 845 1246 849
rect 1330 845 1364 849
rect 1421 808 1455 1090
rect 1512 1049 1546 1053
rect 1630 1049 1664 1053
rect 1506 1037 1552 1049
rect 1506 861 1512 1037
rect 1546 861 1552 1037
rect 1506 849 1552 861
rect 1624 1037 1670 1049
rect 1624 861 1630 1037
rect 1664 861 1670 1037
rect 1624 849 1670 861
rect 1512 845 1546 849
rect 1630 845 1664 849
rect 1721 808 1755 1090
rect 1812 1049 1846 1053
rect 1930 1049 1964 1053
rect 1806 1037 1852 1049
rect 1806 861 1812 1037
rect 1846 861 1852 1037
rect 1806 849 1852 861
rect 1924 1037 1970 1049
rect 1924 861 1930 1037
rect 1964 861 1970 1037
rect 1924 849 1970 861
rect 1812 845 1846 849
rect 1930 845 1964 849
rect 2021 808 2055 1090
rect 2112 1049 2146 1053
rect 2230 1049 2264 1053
rect 2106 1037 2152 1049
rect 2106 861 2112 1037
rect 2146 861 2152 1037
rect 2106 849 2152 861
rect 2224 1037 2270 1049
rect 2224 861 2230 1037
rect 2264 861 2270 1037
rect 2224 849 2270 861
rect 2112 845 2146 849
rect 2230 845 2264 849
rect 2321 808 2355 1090
rect 2412 1049 2446 1053
rect 2406 1037 2452 1049
rect 2406 861 2412 1037
rect 2446 861 2452 1037
rect 2406 849 2452 861
rect 2412 845 2446 849
rect 192 802 284 808
rect 192 768 204 802
rect 272 768 284 802
rect 192 762 284 768
rect 492 802 584 808
rect 492 768 504 802
rect 572 768 584 802
rect 492 762 584 768
rect 792 802 884 808
rect 792 768 804 802
rect 872 768 884 802
rect 792 762 884 768
rect 1092 802 1184 808
rect 1092 768 1104 802
rect 1172 768 1184 802
rect 1092 762 1184 768
rect 1392 802 1484 808
rect 1392 768 1404 802
rect 1472 768 1484 802
rect 1392 762 1484 768
rect 1692 802 1784 808
rect 1692 768 1704 802
rect 1772 768 1784 802
rect 1692 762 1784 768
rect 1992 802 2084 808
rect 1992 768 2004 802
rect 2072 768 2084 802
rect 1992 762 2084 768
rect 2292 802 2384 808
rect 2292 768 2304 802
rect 2372 768 2384 802
rect 2292 762 2384 768
rect 192 415 284 421
rect 192 381 204 415
rect 272 381 284 415
rect 192 375 284 381
rect 492 415 584 421
rect 492 381 504 415
rect 572 381 584 415
rect 492 375 584 381
rect 792 415 884 421
rect 792 381 804 415
rect 872 381 884 415
rect 792 375 884 381
rect 1092 415 1184 421
rect 1092 381 1104 415
rect 1172 381 1184 415
rect 1092 375 1184 381
rect 1392 415 1484 421
rect 1392 381 1404 415
rect 1472 381 1484 415
rect 1392 375 1484 381
rect 1692 415 1784 421
rect 1692 381 1704 415
rect 1772 381 1784 415
rect 1692 375 1784 381
rect 1992 415 2084 421
rect 1992 381 2004 415
rect 2072 381 2084 415
rect 1992 375 2084 381
rect 2292 415 2384 421
rect 2292 381 2304 415
rect 2372 381 2384 415
rect 2292 375 2384 381
rect 130 343 164 347
rect 124 331 170 343
rect 124 225 130 331
rect 164 225 170 331
rect 124 213 170 225
rect 130 209 164 213
rect 221 181 255 375
rect 312 343 346 347
rect 430 343 464 347
rect 306 331 352 343
rect 306 225 312 331
rect 346 225 352 331
rect 306 213 352 225
rect 424 331 470 343
rect 424 225 430 331
rect 464 225 470 331
rect 424 213 470 225
rect 312 209 346 213
rect 430 209 464 213
rect 521 181 555 375
rect 612 343 646 347
rect 730 343 764 347
rect 606 331 652 343
rect 606 225 612 331
rect 646 225 652 331
rect 606 213 652 225
rect 724 331 770 343
rect 724 225 730 331
rect 764 225 770 331
rect 724 213 770 225
rect 612 209 646 213
rect 730 209 764 213
rect 821 181 855 375
rect 912 343 946 347
rect 1030 343 1064 347
rect 906 331 952 343
rect 906 225 912 331
rect 946 225 952 331
rect 906 213 952 225
rect 1024 331 1070 343
rect 1024 225 1030 331
rect 1064 225 1070 331
rect 1024 213 1070 225
rect 912 209 946 213
rect 1030 209 1064 213
rect 1121 181 1155 375
rect 1212 343 1246 347
rect 1330 343 1364 347
rect 1206 331 1252 343
rect 1206 225 1212 331
rect 1246 225 1252 331
rect 1206 213 1252 225
rect 1324 331 1370 343
rect 1324 225 1330 331
rect 1364 225 1370 331
rect 1324 213 1370 225
rect 1212 209 1246 213
rect 1330 209 1364 213
rect 1421 181 1455 375
rect 1512 343 1546 347
rect 1630 343 1664 347
rect 1506 331 1552 343
rect 1506 225 1512 331
rect 1546 225 1552 331
rect 1506 213 1552 225
rect 1624 331 1670 343
rect 1624 225 1630 331
rect 1664 225 1670 331
rect 1624 213 1670 225
rect 1512 209 1546 213
rect 1630 209 1664 213
rect 1721 181 1755 375
rect 1812 343 1846 347
rect 1930 343 1964 347
rect 1806 331 1852 343
rect 1806 225 1812 331
rect 1846 225 1852 331
rect 1806 213 1852 225
rect 1924 331 1970 343
rect 1924 225 1930 331
rect 1964 225 1970 331
rect 1924 213 1970 225
rect 1812 209 1846 213
rect 1930 209 1964 213
rect 2021 181 2055 375
rect 2112 343 2146 347
rect 2230 343 2264 347
rect 2106 331 2152 343
rect 2106 225 2112 331
rect 2146 225 2152 331
rect 2106 213 2152 225
rect 2224 331 2270 343
rect 2224 225 2230 331
rect 2264 225 2270 331
rect 2224 213 2270 225
rect 2112 209 2146 213
rect 2230 209 2264 213
rect 2321 181 2355 375
rect 2412 343 2446 347
rect 2406 331 2452 343
rect 2406 225 2412 331
rect 2446 225 2452 331
rect 2406 213 2452 225
rect 2412 209 2446 213
rect 192 175 284 181
rect 192 141 204 175
rect 272 141 284 175
rect 192 135 284 141
rect 492 175 584 181
rect 492 141 504 175
rect 572 141 584 175
rect 492 135 584 141
rect 792 175 884 181
rect 792 141 804 175
rect 872 141 884 175
rect 792 135 884 141
rect 1092 175 1184 181
rect 1092 141 1104 175
rect 1172 141 1184 175
rect 1092 135 1184 141
rect 1392 175 1484 181
rect 1392 141 1404 175
rect 1472 141 1484 175
rect 1392 135 1484 141
rect 1692 175 1784 181
rect 1692 141 1704 175
rect 1772 141 1784 175
rect 1692 135 1784 141
rect 1992 175 2084 181
rect 1992 141 2004 175
rect 2072 141 2084 175
rect 1992 135 2084 141
rect 2292 175 2384 181
rect 2292 141 2304 175
rect 2372 141 2384 175
rect 2292 135 2384 141
rect 88 82 2488 94
rect 88 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2488 82
rect 88 36 2488 48
<< labels >>
flabel metal1 88 1168 2488 1226 0 FreeSans 256 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal1 88 36 2488 94 0 FreeSans 256 0 0 0 VSS
port 1 nsew ground bidirectional
<< end >>
