magic
tech sky130A
magscale 1 2
timestamp 1727641773
<< dnwell >>
rect -606 -335 3302 1898
<< nwell >>
rect -686 1692 3382 1978
rect -686 -129 -400 1692
rect 3096 -129 3382 1692
rect -686 -415 3382 -129
<< nsubdiff >>
rect -649 1921 3345 1941
rect -649 1887 -569 1921
rect 3265 1887 3345 1921
rect -649 1867 3345 1887
rect -649 1861 -575 1867
rect -649 -298 -629 1861
rect -595 -298 -575 1861
rect -649 -304 -575 -298
rect 3271 1861 3345 1867
rect 3271 -298 3291 1861
rect 3325 -298 3345 1861
rect 3271 -304 3345 -298
rect -649 -324 3345 -304
rect -649 -358 -569 -324
rect 3265 -358 3345 -324
rect -649 -378 3345 -358
<< nsubdiffcont >>
rect -569 1887 3265 1921
rect -629 -298 -595 1861
rect 3291 -298 3325 1861
rect -569 -358 3265 -324
<< locali >>
rect -629 1887 -569 1921
rect 3265 1887 3325 1921
rect -629 1861 -595 1887
rect -629 -324 -595 -298
rect 3291 1861 3325 1887
rect 3291 -324 3325 -298
rect -629 -358 -569 -324
rect 3265 -358 3325 -324
use tie_highs  tie_highs_0
timestamp 1727641773
transform 1 0 60 0 1 0
box -60 0 2636 1292
<< end >>
