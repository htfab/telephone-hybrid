magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< metal1 >>
rect 0 44952 200 45152
rect 28872 44952 29072 45152
rect 7861 41394 7867 41446
rect 7919 41394 7925 41446
rect 8161 41394 8167 41446
rect 8219 41394 8225 41446
rect 8461 41394 8467 41446
rect 8519 41394 8525 41446
rect 8761 41394 8767 41446
rect 8819 41394 8825 41446
rect 9061 41394 9067 41446
rect 9119 41394 9125 41446
rect 9361 41394 9367 41446
rect 9419 41394 9425 41446
rect 9661 41394 9667 41446
rect 9719 41394 9725 41446
rect 9961 41394 9967 41446
rect 10019 41394 10025 41446
rect 13061 41394 13067 41446
rect 13119 41394 13125 41446
rect 13361 41394 13367 41446
rect 13419 41394 13425 41446
rect 13661 41394 13667 41446
rect 13719 41394 13725 41446
rect 13961 41394 13967 41446
rect 14019 41394 14025 41446
rect 14261 41394 14267 41446
rect 14319 41394 14325 41446
rect 14561 41394 14567 41446
rect 14619 41394 14625 41446
rect 14861 41394 14867 41446
rect 14919 41394 14925 41446
rect 15161 41394 15167 41446
rect 15219 41394 15225 41446
rect 2834 41100 2840 41170
rect 2910 41100 2916 41170
rect 3134 41100 3140 41170
rect 3210 41100 3216 41170
rect 3434 41100 3440 41170
rect 3510 41100 3516 41170
rect 3734 41100 3740 41170
rect 3810 41100 3816 41170
rect 4034 41100 4040 41170
rect 4110 41100 4116 41170
rect 4334 41100 4340 41170
rect 4410 41100 4416 41170
rect 4634 41100 4640 41170
rect 4710 41100 4716 41170
rect 4934 41100 4940 41170
rect 5010 41100 5016 41170
rect 21552 41161 21558 41213
rect 21610 41161 21616 41213
rect 21852 41161 21858 41213
rect 21910 41161 21916 41213
rect 22152 41161 22158 41213
rect 22210 41161 22216 41213
rect 22452 41161 22458 41213
rect 22510 41161 22516 41213
rect 22752 41161 22758 41213
rect 22810 41161 22816 41213
rect 23052 41161 23058 41213
rect 23110 41161 23116 41213
rect 23352 41161 23358 41213
rect 23410 41161 23416 41213
rect 23652 41161 23658 41213
rect 23710 41161 23716 41213
rect 7958 35757 8010 35763
rect 7958 35699 8010 35705
rect 8258 35757 8310 35763
rect 8258 35699 8310 35705
rect 8558 35757 8610 35763
rect 8558 35699 8610 35705
rect 8858 35757 8910 35763
rect 8858 35699 8910 35705
rect 9158 35757 9210 35763
rect 9158 35699 9210 35705
rect 9458 35757 9510 35763
rect 9458 35699 9510 35705
rect 9758 35757 9810 35763
rect 9758 35699 9810 35705
rect 10058 35757 10110 35763
rect 10058 35699 10110 35705
rect 13158 35757 13210 35763
rect 13158 35699 13210 35705
rect 13458 35757 13510 35763
rect 13458 35699 13510 35705
rect 13758 35757 13810 35763
rect 13758 35699 13810 35705
rect 14058 35757 14110 35763
rect 14058 35699 14110 35705
rect 14358 35757 14410 35763
rect 14358 35699 14410 35705
rect 14658 35757 14710 35763
rect 14658 35699 14710 35705
rect 14958 35757 15010 35763
rect 14958 35699 15010 35705
rect 15258 35757 15310 35763
rect 15258 35699 15310 35705
rect 21658 35538 21692 35635
rect 21958 35538 21992 35635
rect 22258 35538 22292 35635
rect 22558 35538 22592 35635
rect 22858 35538 22892 35635
rect 23158 35538 23192 35635
rect 23458 35538 23492 35635
rect 23758 35538 23792 35635
rect 21649 35532 21701 35538
rect 21649 35474 21701 35480
rect 21949 35532 22001 35538
rect 21949 35474 22001 35480
rect 22249 35532 22301 35538
rect 22249 35474 22301 35480
rect 22549 35532 22601 35538
rect 22549 35474 22601 35480
rect 22849 35532 22901 35538
rect 22849 35474 22901 35480
rect 23149 35532 23201 35538
rect 23149 35474 23201 35480
rect 23449 35532 23501 35538
rect 23449 35474 23501 35480
rect 23749 35532 23801 35538
rect 23749 35474 23801 35480
rect 7719 33569 7789 33575
rect 8631 33569 8701 33575
rect 7789 33499 8631 33569
rect 7719 33493 7789 33499
rect 8631 33493 8701 33499
rect 8175 33369 8245 33375
rect 13999 33369 14069 33375
rect 8245 33299 13999 33369
rect 8175 33293 8245 33299
rect 13999 33293 14069 33299
rect 7934 33169 8004 33175
rect 8390 33169 8460 33175
rect 8004 33099 8390 33169
rect 7934 33093 8004 33099
rect 8390 33093 8460 33099
rect 8846 32969 8916 32975
rect 13302 32969 13372 32975
rect 8916 32899 13302 32969
rect 8846 32893 8916 32899
rect 13302 32893 13372 32899
rect 9061 32769 9131 32775
rect 9973 32769 10043 32775
rect 9131 32699 9973 32769
rect 9061 32693 9131 32699
rect 9973 32693 10043 32699
rect 9517 32569 9587 32575
rect 15341 32569 15411 32575
rect 9587 32499 15341 32569
rect 9517 32493 9587 32499
rect 15341 32493 15411 32499
rect 9276 32369 9346 32375
rect 9732 32369 9802 32375
rect 9346 32299 9732 32369
rect 9276 32293 9346 32299
rect 9732 32293 9802 32299
rect 10188 32169 10258 32175
rect 14644 32169 14714 32175
rect 10258 32099 14644 32169
rect 10188 32093 10258 32099
rect 14644 32093 14714 32099
rect 5947 31969 6017 31975
rect 13087 31969 13157 31975
rect 6017 31899 13087 31969
rect 5947 31893 6017 31899
rect 13087 31893 13157 31899
rect 11315 31769 11385 31775
rect 13543 31769 13613 31775
rect 11385 31699 13543 31769
rect 11315 31693 11385 31699
rect 13543 31693 13613 31699
rect 5250 31569 5320 31575
rect 13758 31569 13828 31575
rect 5320 31499 13758 31569
rect 5250 31493 5320 31499
rect 13758 31493 13828 31499
rect 10618 31369 10688 31375
rect 14214 31369 14284 31375
rect 10688 31299 14214 31369
rect 10618 31293 10688 31299
rect 14214 31293 14284 31299
rect 7289 31169 7359 31175
rect 14429 31169 14499 31175
rect 7359 31099 14429 31169
rect 7289 31093 7359 31099
rect 14429 31093 14499 31099
rect 12657 30969 12727 30975
rect 14885 30969 14955 30975
rect 12727 30899 14885 30969
rect 12657 30893 12727 30899
rect 14885 30893 14955 30899
rect 6592 30769 6662 30775
rect 15100 30769 15170 30775
rect 6662 30699 15100 30769
rect 6592 30693 6662 30699
rect 15100 30693 15170 30699
rect 11960 30569 12030 30575
rect 15556 30569 15626 30575
rect 12030 30499 15556 30569
rect 11960 30493 12030 30499
rect 15556 30493 15626 30499
rect 18025 25029 18095 25035
rect 18095 24959 21640 25029
rect 21710 24959 21716 25029
rect 18025 24953 18095 24959
rect 13999 24729 14069 24735
rect 14069 24659 21940 24729
rect 22010 24659 22016 24729
rect 13999 24653 14069 24659
rect 15341 24429 15411 24435
rect 15411 24359 22240 24429
rect 22310 24359 22316 24429
rect 15341 24353 15411 24359
rect 16683 24129 16753 24135
rect 16936 24129 17006 24135
rect 16753 24059 16936 24129
rect 17006 24059 22540 24129
rect 22610 24059 22616 24129
rect 16683 24053 16753 24059
rect 16936 24053 17006 24059
rect 3202 23829 3272 23835
rect 3272 23759 22840 23829
rect 22910 23759 22916 23829
rect 3202 23753 3272 23759
rect 3502 23529 3572 23535
rect 3572 23459 23140 23529
rect 23210 23459 23216 23529
rect 3502 23453 3572 23459
rect 3802 23229 3872 23235
rect 3872 23159 23440 23229
rect 23510 23159 23516 23229
rect 3802 23153 3872 23159
rect 4102 22929 4172 22935
rect 4172 22859 23740 22929
rect 23810 22859 23816 22929
rect 4102 22853 4172 22859
rect 3502 11515 3572 11521
rect 3572 11506 5936 11515
rect 3572 11454 5875 11506
rect 5927 11454 5936 11506
rect 3572 11445 5936 11454
rect 3502 11439 3572 11445
rect 3802 10173 3872 10179
rect 3872 10164 5936 10173
rect 3872 10112 5875 10164
rect 5927 10112 5936 10164
rect 3872 10103 5936 10112
rect 3802 10097 3872 10103
rect 12428 9916 12434 10016
rect 12534 9916 12540 10016
rect 4102 8831 4172 8837
rect 4172 8822 5936 8831
rect 4172 8770 5875 8822
rect 5927 8770 5936 8822
rect 4172 8761 5936 8770
rect 4102 8755 4172 8761
rect 3201 7489 3271 7495
rect 3271 7480 5936 7489
rect 3271 7428 5875 7480
rect 5927 7428 5936 7480
rect 3271 7419 5936 7428
rect 3201 7413 3271 7419
rect 0 0 200 200
rect 28872 0 29072 200
<< via1 >>
rect 7867 41394 7919 41446
rect 8167 41394 8219 41446
rect 8467 41394 8519 41446
rect 8767 41394 8819 41446
rect 9067 41394 9119 41446
rect 9367 41394 9419 41446
rect 9667 41394 9719 41446
rect 9967 41394 10019 41446
rect 13067 41394 13119 41446
rect 13367 41394 13419 41446
rect 13667 41394 13719 41446
rect 13967 41394 14019 41446
rect 14267 41394 14319 41446
rect 14567 41394 14619 41446
rect 14867 41394 14919 41446
rect 15167 41394 15219 41446
rect 2840 41100 2910 41170
rect 3140 41100 3210 41170
rect 3440 41100 3510 41170
rect 3740 41100 3810 41170
rect 4040 41100 4110 41170
rect 4340 41100 4410 41170
rect 4640 41100 4710 41170
rect 4940 41100 5010 41170
rect 21558 41161 21610 41213
rect 21858 41161 21910 41213
rect 22158 41161 22210 41213
rect 22458 41161 22510 41213
rect 22758 41161 22810 41213
rect 23058 41161 23110 41213
rect 23358 41161 23410 41213
rect 23658 41161 23710 41213
rect 7958 35705 8010 35757
rect 8258 35705 8310 35757
rect 8558 35705 8610 35757
rect 8858 35705 8910 35757
rect 9158 35705 9210 35757
rect 9458 35705 9510 35757
rect 9758 35705 9810 35757
rect 10058 35705 10110 35757
rect 13158 35705 13210 35757
rect 13458 35705 13510 35757
rect 13758 35705 13810 35757
rect 14058 35705 14110 35757
rect 14358 35705 14410 35757
rect 14658 35705 14710 35757
rect 14958 35705 15010 35757
rect 15258 35705 15310 35757
rect 21649 35480 21701 35532
rect 21949 35480 22001 35532
rect 22249 35480 22301 35532
rect 22549 35480 22601 35532
rect 22849 35480 22901 35532
rect 23149 35480 23201 35532
rect 23449 35480 23501 35532
rect 23749 35480 23801 35532
rect 7719 33499 7789 33569
rect 8631 33499 8701 33569
rect 8175 33299 8245 33369
rect 13999 33299 14069 33369
rect 7934 33099 8004 33169
rect 8390 33099 8460 33169
rect 8846 32899 8916 32969
rect 13302 32899 13372 32969
rect 9061 32699 9131 32769
rect 9973 32699 10043 32769
rect 9517 32499 9587 32569
rect 15341 32499 15411 32569
rect 9276 32299 9346 32369
rect 9732 32299 9802 32369
rect 10188 32099 10258 32169
rect 14644 32099 14714 32169
rect 5947 31899 6017 31969
rect 13087 31899 13157 31969
rect 11315 31699 11385 31769
rect 13543 31699 13613 31769
rect 5250 31499 5320 31569
rect 13758 31499 13828 31569
rect 10618 31299 10688 31369
rect 14214 31299 14284 31369
rect 7289 31099 7359 31169
rect 14429 31099 14499 31169
rect 12657 30899 12727 30969
rect 14885 30899 14955 30969
rect 6592 30699 6662 30769
rect 15100 30699 15170 30769
rect 11960 30499 12030 30569
rect 15556 30499 15626 30569
rect 18025 24959 18095 25029
rect 21640 24959 21710 25029
rect 13999 24659 14069 24729
rect 21940 24659 22010 24729
rect 15341 24359 15411 24429
rect 22240 24359 22310 24429
rect 16683 24059 16753 24129
rect 16936 24059 17006 24129
rect 22540 24059 22610 24129
rect 3202 23759 3272 23829
rect 22840 23759 22910 23829
rect 3502 23459 3572 23529
rect 23140 23459 23210 23529
rect 3802 23159 3872 23229
rect 23440 23159 23510 23229
rect 4102 22859 4172 22929
rect 23740 22859 23810 22929
rect 3502 11445 3572 11515
rect 5875 11454 5927 11506
rect 3802 10103 3872 10173
rect 5875 10112 5927 10164
rect 12434 9916 12534 10016
rect 4102 8761 4172 8831
rect 5875 8770 5927 8822
rect 3201 7419 3271 7489
rect 5875 7428 5927 7480
<< metal2 >>
rect 3001 44674 3071 44679
rect 3553 44674 3623 44679
rect 4105 44674 4175 44679
rect 4657 44674 4727 44679
rect 5209 44674 5279 44679
rect 5761 44674 5831 44679
rect 6313 44674 6383 44679
rect 6865 44674 6935 44679
rect 7417 44674 7487 44679
rect 7969 44674 8039 44679
rect 8521 44674 8591 44679
rect 9073 44674 9143 44679
rect 9625 44674 9695 44679
rect 10177 44674 10247 44679
rect 10729 44674 10799 44679
rect 11281 44674 11351 44679
rect 11833 44674 11903 44679
rect 12385 44674 12455 44679
rect 12937 44674 13007 44679
rect 13489 44674 13559 44679
rect 14041 44674 14111 44679
rect 14593 44674 14663 44679
rect 15145 44674 15215 44679
rect 15697 44674 15767 44679
rect 20665 44674 20735 44679
rect 21217 44674 21287 44679
rect 21769 44674 21839 44679
rect 22321 44674 22391 44679
rect 22873 44674 22943 44679
rect 23425 44674 23495 44679
rect 23977 44674 24047 44679
rect 24529 44674 24599 44679
rect 2997 44614 3006 44674
rect 3066 44614 3075 44674
rect 3549 44614 3558 44674
rect 3618 44614 3627 44674
rect 4101 44614 4110 44674
rect 4170 44614 4179 44674
rect 4653 44614 4662 44674
rect 4722 44614 4731 44674
rect 5205 44614 5214 44674
rect 5274 44614 5283 44674
rect 5757 44614 5766 44674
rect 5826 44614 5835 44674
rect 6309 44614 6318 44674
rect 6378 44614 6387 44674
rect 6861 44614 6870 44674
rect 6930 44614 6939 44674
rect 7413 44614 7422 44674
rect 7482 44614 7491 44674
rect 7965 44614 7974 44674
rect 8034 44614 8043 44674
rect 8517 44614 8526 44674
rect 8586 44614 8595 44674
rect 9069 44614 9078 44674
rect 9138 44614 9147 44674
rect 9621 44614 9630 44674
rect 9690 44614 9699 44674
rect 10173 44614 10182 44674
rect 10242 44614 10251 44674
rect 10725 44614 10734 44674
rect 10794 44614 10803 44674
rect 11277 44614 11286 44674
rect 11346 44614 11355 44674
rect 11829 44614 11838 44674
rect 11898 44614 11907 44674
rect 12381 44614 12390 44674
rect 12450 44614 12459 44674
rect 12933 44614 12942 44674
rect 13002 44614 13011 44674
rect 13485 44614 13494 44674
rect 13554 44614 13563 44674
rect 14037 44614 14046 44674
rect 14106 44614 14115 44674
rect 14589 44614 14598 44674
rect 14658 44614 14667 44674
rect 15141 44614 15150 44674
rect 15210 44614 15219 44674
rect 15693 44614 15702 44674
rect 15762 44614 15771 44674
rect 20661 44614 20670 44674
rect 20730 44614 20739 44674
rect 21213 44614 21222 44674
rect 21282 44614 21291 44674
rect 21765 44614 21774 44674
rect 21834 44614 21843 44674
rect 22317 44614 22326 44674
rect 22386 44614 22395 44674
rect 22869 44614 22878 44674
rect 22938 44614 22947 44674
rect 23421 44614 23430 44674
rect 23490 44614 23499 44674
rect 23973 44614 23982 44674
rect 24042 44614 24051 44674
rect 24525 44614 24534 44674
rect 24594 44614 24603 44674
rect 3001 44082 3071 44614
rect 3000 43741 3071 44082
rect 2840 43671 3071 43741
rect 2840 41170 2910 43671
rect 3553 43541 3623 44614
rect 2840 41094 2910 41100
rect 3140 43471 3623 43541
rect 3140 41170 3210 43471
rect 4105 43341 4175 44614
rect 3140 41094 3210 41100
rect 3440 43271 4175 43341
rect 3440 41170 3510 43271
rect 4657 43141 4727 44614
rect 3440 41094 3510 41100
rect 3740 43071 4727 43141
rect 3740 41170 3810 43071
rect 5209 42941 5279 44614
rect 3740 41094 3810 41100
rect 4040 42871 5279 42941
rect 4040 41170 4110 42871
rect 5761 42741 5831 44614
rect 4040 41094 4110 41100
rect 4340 42671 5831 42741
rect 4340 41170 4410 42671
rect 6313 42541 6383 44614
rect 4340 41094 4410 41100
rect 4640 42471 6383 42541
rect 4640 41170 4710 42471
rect 6865 42341 6935 44614
rect 4640 41094 4710 41100
rect 4940 42271 6935 42341
rect 7417 42341 7487 44614
rect 7969 42541 8039 44614
rect 8521 43341 8591 44614
rect 8458 43271 8591 43341
rect 7969 42473 8228 42541
rect 8008 42471 8228 42473
rect 7417 42271 7928 42341
rect 4940 41170 5010 42271
rect 7858 41446 7928 42271
rect 7858 41394 7867 41446
rect 7919 41394 7928 41446
rect 7858 41385 7928 41394
rect 8158 41446 8228 42471
rect 8158 41394 8167 41446
rect 8219 41394 8228 41446
rect 8158 41385 8228 41394
rect 8458 41446 8528 43271
rect 9073 43141 9143 44614
rect 8458 41394 8467 41446
rect 8519 41394 8528 41446
rect 8458 41385 8528 41394
rect 8758 43071 9143 43141
rect 8758 41446 8828 43071
rect 9625 42941 9695 44614
rect 8758 41394 8767 41446
rect 8819 41394 8828 41446
rect 8758 41385 8828 41394
rect 9058 42871 9695 42941
rect 9058 41446 9128 42871
rect 10177 42741 10247 44614
rect 9058 41394 9067 41446
rect 9119 41394 9128 41446
rect 9058 41385 9128 41394
rect 9358 42671 10247 42741
rect 9358 41446 9428 42671
rect 10729 42541 10799 44614
rect 9358 41394 9367 41446
rect 9419 41394 9428 41446
rect 9358 41385 9428 41394
rect 9658 42471 10799 42541
rect 9658 41446 9728 42471
rect 11281 42341 11351 44614
rect 9658 41394 9667 41446
rect 9719 41394 9728 41446
rect 9658 41385 9728 41394
rect 9958 42271 11351 42341
rect 11833 42341 11903 44614
rect 12385 42541 12455 44614
rect 12937 42741 13007 44614
rect 13489 42941 13559 44614
rect 14041 43141 14111 44614
rect 14041 43071 14328 43141
rect 13489 42871 14028 42941
rect 12937 42671 13728 42741
rect 12385 42471 13428 42541
rect 11833 42271 13128 42341
rect 9958 41446 10028 42271
rect 9958 41394 9967 41446
rect 10019 41394 10028 41446
rect 9958 41385 10028 41394
rect 13058 41446 13128 42271
rect 13058 41394 13067 41446
rect 13119 41394 13128 41446
rect 13058 41385 13128 41394
rect 13358 41446 13428 42471
rect 13358 41394 13367 41446
rect 13419 41394 13428 41446
rect 13358 41385 13428 41394
rect 13658 41446 13728 42671
rect 13658 41394 13667 41446
rect 13719 41394 13728 41446
rect 13658 41385 13728 41394
rect 13958 41446 14028 42871
rect 13958 41394 13967 41446
rect 14019 41394 14028 41446
rect 13958 41385 14028 41394
rect 14258 41446 14328 43071
rect 14593 42741 14663 44614
rect 14258 41394 14267 41446
rect 14319 41394 14328 41446
rect 14258 41385 14328 41394
rect 14558 42671 14663 42741
rect 14558 41446 14628 42671
rect 15145 42541 15215 44614
rect 14558 41394 14567 41446
rect 14619 41394 14628 41446
rect 14558 41385 14628 41394
rect 14858 42471 15215 42541
rect 14858 41446 14928 42471
rect 14858 41394 14867 41446
rect 14919 41394 14928 41446
rect 14858 41385 14928 41394
rect 15158 42340 15228 42341
rect 15697 42340 15767 44614
rect 15158 42271 15767 42340
rect 20665 42341 20735 44614
rect 21217 42541 21287 44614
rect 21769 42741 21839 44614
rect 22321 42941 22391 44614
rect 22873 42941 22943 44614
rect 22321 42871 22519 42941
rect 21769 42671 22219 42741
rect 21217 42471 21919 42541
rect 20665 42271 21619 42341
rect 15158 42270 15728 42271
rect 15158 41446 15228 42270
rect 15158 41394 15167 41446
rect 15219 41394 15228 41446
rect 15158 41385 15228 41394
rect 21549 41227 21619 42271
rect 21849 41227 21919 42471
rect 22149 41227 22219 42671
rect 22449 41227 22519 42871
rect 22749 42871 22943 42941
rect 22749 41227 22819 42871
rect 23425 42741 23495 44614
rect 23049 42671 23495 42741
rect 23049 41227 23119 42671
rect 23977 42541 24047 44614
rect 23349 42471 24047 42541
rect 23349 41227 23419 42471
rect 24529 42341 24599 44614
rect 23649 42271 24599 42341
rect 23649 41227 23719 42271
rect 21544 41213 21624 41227
rect 21544 41161 21558 41213
rect 21610 41161 21624 41213
rect 21544 41147 21624 41161
rect 21844 41213 21924 41227
rect 21844 41161 21858 41213
rect 21910 41161 21924 41213
rect 21844 41147 21924 41161
rect 22144 41213 22224 41227
rect 22144 41161 22158 41213
rect 22210 41161 22224 41213
rect 22144 41147 22224 41161
rect 22444 41213 22524 41227
rect 22444 41161 22458 41213
rect 22510 41161 22524 41213
rect 22444 41147 22524 41161
rect 22744 41213 22824 41227
rect 22744 41161 22758 41213
rect 22810 41161 22824 41213
rect 22744 41147 22824 41161
rect 23044 41213 23124 41227
rect 23044 41161 23058 41213
rect 23110 41161 23124 41213
rect 23044 41147 23124 41161
rect 23344 41213 23424 41227
rect 23344 41161 23358 41213
rect 23410 41161 23424 41213
rect 23344 41147 23424 41161
rect 23644 41213 23724 41227
rect 23644 41161 23658 41213
rect 23710 41161 23724 41213
rect 23644 41147 23724 41161
rect 4940 41094 5010 41100
rect 7949 35757 8019 35766
rect 7949 35705 7958 35757
rect 8010 35705 8019 35757
rect 7949 34369 8019 35705
rect 7719 34299 8019 34369
rect 8249 35757 8319 35766
rect 8249 35705 8258 35757
rect 8310 35705 8319 35757
rect 7719 33569 7789 34299
rect 8249 34169 8319 35705
rect 8175 34099 8319 34169
rect 8549 35757 8619 35766
rect 8549 35705 8558 35757
rect 8610 35705 8619 35757
rect 7713 33499 7719 33569
rect 7789 33499 7795 33569
rect 8175 33369 8245 34099
rect 8549 33969 8619 35705
rect 8849 35757 8919 35766
rect 8849 35705 8858 35757
rect 8910 35705 8919 35757
rect 8849 33969 8919 35705
rect 9149 35757 9219 35766
rect 9149 35705 9158 35757
rect 9210 35705 9219 35757
rect 9149 33969 9219 35705
rect 8390 33899 8619 33969
rect 8846 33899 8919 33969
rect 9061 33899 9219 33969
rect 9449 35757 9519 35766
rect 9449 35705 9458 35757
rect 9510 35705 9519 35757
rect 9449 33969 9519 35705
rect 9749 35757 9819 35766
rect 9749 35705 9758 35757
rect 9810 35705 9819 35757
rect 9749 33969 9819 35705
rect 9449 33899 9587 33969
rect 8169 33299 8175 33369
rect 8245 33299 8251 33369
rect 8390 33169 8460 33899
rect 8625 33499 8631 33569
rect 8701 33499 8707 33569
rect 7928 33099 7934 33169
rect 8004 33099 8010 33169
rect 8384 33099 8390 33169
rect 8460 33099 8466 33169
rect 5941 31899 5947 31969
rect 6017 31899 6023 31969
rect 5244 31499 5250 31569
rect 5320 31499 5326 31569
rect 5250 29627 5320 31499
rect 5947 29627 6017 31899
rect 7283 31099 7289 31169
rect 7359 31099 7365 31169
rect 6586 30699 6592 30769
rect 6662 30699 6668 30769
rect 6592 29627 6662 30699
rect 7289 29627 7359 31099
rect 7934 29627 8004 33099
rect 8631 29627 8701 33499
rect 8846 32969 8916 33899
rect 8840 32899 8846 32969
rect 8916 32899 8922 32969
rect 9061 32769 9131 33899
rect 9055 32699 9061 32769
rect 9131 32699 9137 32769
rect 9517 32569 9587 33899
rect 9732 33899 9819 33969
rect 10049 35757 10119 35766
rect 10049 35705 10058 35757
rect 10110 35705 10119 35757
rect 10049 33969 10119 35705
rect 13149 35757 13219 35766
rect 13149 35705 13158 35757
rect 13210 35705 13219 35757
rect 13149 33969 13219 35705
rect 10049 33899 10258 33969
rect 9511 32499 9517 32569
rect 9587 32499 9593 32569
rect 9732 32369 9802 33899
rect 9967 32699 9973 32769
rect 10043 32699 10049 32769
rect 9270 32299 9276 32369
rect 9346 32299 9352 32369
rect 9726 32299 9732 32369
rect 9802 32299 9808 32369
rect 9276 29627 9346 32299
rect 9973 29627 10043 32699
rect 10188 32169 10258 33899
rect 13087 33899 13219 33969
rect 13449 35757 13519 35766
rect 13449 35705 13458 35757
rect 13510 35705 13519 35757
rect 13449 33969 13519 35705
rect 13749 35757 13819 35766
rect 13749 35705 13758 35757
rect 13810 35705 13819 35757
rect 13749 33969 13819 35705
rect 14049 35757 14119 35766
rect 14049 35705 14058 35757
rect 14110 35705 14119 35757
rect 14049 33969 14119 35705
rect 14349 35757 14419 35766
rect 14349 35705 14358 35757
rect 14410 35705 14419 35757
rect 14349 34169 14419 35705
rect 14649 35757 14719 35766
rect 14649 35705 14658 35757
rect 14710 35705 14719 35757
rect 14349 34099 14499 34169
rect 13449 33899 13613 33969
rect 13749 33899 13828 33969
rect 14049 33899 14284 33969
rect 10182 32099 10188 32169
rect 10258 32099 10264 32169
rect 13087 31969 13157 33899
rect 13296 32899 13302 32969
rect 13372 32899 13378 32969
rect 13081 31899 13087 31969
rect 13157 31899 13163 31969
rect 11309 31699 11315 31769
rect 11385 31699 11391 31769
rect 10612 31299 10618 31369
rect 10688 31299 10694 31369
rect 10618 29627 10688 31299
rect 11315 29627 11385 31699
rect 12651 30899 12657 30969
rect 12727 30899 12733 30969
rect 11954 30499 11960 30569
rect 12030 30499 12036 30569
rect 11960 29627 12030 30499
rect 12657 29627 12727 30899
rect 13302 29627 13372 32899
rect 13543 31769 13613 33899
rect 13537 31699 13543 31769
rect 13613 31699 13619 31769
rect 13758 31569 13828 33899
rect 13993 33299 13999 33369
rect 14069 33299 14075 33369
rect 13752 31499 13758 31569
rect 13828 31499 13834 31569
rect 13999 29627 14069 33299
rect 14214 31369 14284 33899
rect 14208 31299 14214 31369
rect 14284 31299 14290 31369
rect 14429 31169 14499 34099
rect 14649 33969 14719 35705
rect 14949 35757 15019 35766
rect 14949 35705 14958 35757
rect 15010 35705 15019 35757
rect 14949 34169 15019 35705
rect 15249 35757 15319 35766
rect 15249 35705 15258 35757
rect 15310 35705 15319 35757
rect 15249 34369 15319 35705
rect 21640 35532 21710 35541
rect 21640 35480 21649 35532
rect 21701 35480 21710 35532
rect 15249 34299 15626 34369
rect 14949 34099 15170 34169
rect 14649 33899 14955 33969
rect 14638 32099 14644 32169
rect 14714 32099 14720 32169
rect 14423 31099 14429 31169
rect 14499 31099 14505 31169
rect 14644 29627 14714 32099
rect 14885 30969 14955 33899
rect 14879 30899 14885 30969
rect 14955 30899 14961 30969
rect 15100 30769 15170 34099
rect 15335 32499 15341 32569
rect 15411 32499 15417 32569
rect 15094 30699 15100 30769
rect 15170 30699 15176 30769
rect 15341 29627 15411 32499
rect 15556 30569 15626 34299
rect 15550 30499 15556 30569
rect 15626 30499 15632 30569
rect 5268 29419 5302 29627
rect 5965 29419 5999 29627
rect 6610 29419 6644 29627
rect 7307 29419 7341 29627
rect 7952 29419 7986 29627
rect 8649 29419 8683 29627
rect 9294 29419 9328 29627
rect 9991 29419 10025 29627
rect 10636 29419 10670 29627
rect 11333 29419 11367 29627
rect 11978 29419 12012 29627
rect 12675 29419 12709 29627
rect 13320 29419 13354 29627
rect 14017 29419 14051 29627
rect 14662 29419 14696 29627
rect 15359 29418 15393 29627
rect 13999 24729 14069 26284
rect 13993 24659 13999 24729
rect 14069 24659 14075 24729
rect 15341 24429 15411 26298
rect 15335 24359 15341 24429
rect 15411 24359 15417 24429
rect 16683 24129 16753 26282
rect 18025 25029 18095 26287
rect 21640 25029 21710 35480
rect 18019 24959 18025 25029
rect 18095 24959 18101 25029
rect 21640 24950 21710 24959
rect 21940 35532 22010 35541
rect 21940 35480 21949 35532
rect 22001 35480 22010 35532
rect 21940 24729 22010 35480
rect 21940 24650 22010 24659
rect 22240 35532 22310 35541
rect 22240 35480 22249 35532
rect 22301 35480 22310 35532
rect 22240 24429 22310 35480
rect 22240 24350 22310 24359
rect 22540 35532 22610 35541
rect 22540 35480 22549 35532
rect 22601 35480 22610 35532
rect 22540 24129 22610 35480
rect 16677 24059 16683 24129
rect 16753 24059 16759 24129
rect 16930 24059 16936 24129
rect 17006 24059 17012 24129
rect 3196 23759 3202 23829
rect 3272 23759 3278 23829
rect 3202 7489 3272 23759
rect 3496 23459 3502 23529
rect 3572 23459 3578 23529
rect 3502 11515 3572 23459
rect 3796 23159 3802 23229
rect 3872 23159 3878 23229
rect 3496 11445 3502 11515
rect 3572 11445 3578 11515
rect 3802 10173 3872 23159
rect 4096 22859 4102 22929
rect 4172 22859 4178 22929
rect 3796 10103 3802 10173
rect 3872 10103 3878 10173
rect 4102 8831 4172 22859
rect 5869 11454 5875 11506
rect 5927 11497 5933 11506
rect 5927 11463 6415 11497
rect 5927 11454 5933 11463
rect 5869 10112 5875 10164
rect 5927 10155 5933 10164
rect 5927 10121 6415 10155
rect 5927 10112 5933 10121
rect 10261 10077 11191 10177
rect 10261 9773 10361 10077
rect 11091 10016 11191 10077
rect 12434 10016 12534 10022
rect 11091 9916 12434 10016
rect 12434 9910 12534 9916
rect 9866 9673 10361 9773
rect 4096 8761 4102 8831
rect 4172 8761 4178 8831
rect 5869 8770 5875 8822
rect 5927 8813 5933 8822
rect 5927 8779 6415 8813
rect 5927 8770 5933 8779
rect 3195 7419 3201 7489
rect 3271 7419 3277 7489
rect 5869 7428 5875 7480
rect 5927 7471 5933 7480
rect 5927 7437 6415 7471
rect 5927 7428 5933 7437
rect 9866 6687 9966 9673
rect 7952 6587 9966 6687
rect 7952 195 8052 6587
rect 16936 5982 17006 24059
rect 22540 24050 22610 24059
rect 22840 35532 22910 35541
rect 22840 35480 22849 35532
rect 22901 35480 22910 35532
rect 22840 23829 22910 35480
rect 22840 23750 22910 23759
rect 23140 35532 23210 35541
rect 23140 35480 23149 35532
rect 23201 35480 23210 35532
rect 23140 23529 23210 35480
rect 23140 23450 23210 23459
rect 23440 35532 23510 35541
rect 23440 35480 23449 35532
rect 23501 35480 23510 35532
rect 23440 23229 23510 35480
rect 23440 23150 23510 23159
rect 23740 35532 23810 35541
rect 23740 35480 23749 35532
rect 23801 35480 23810 35532
rect 23740 22929 23810 35480
rect 23740 22850 23810 22859
rect 21677 8277 27374 8377
rect 21677 7956 21777 8277
rect 16936 5912 17356 5982
rect 16919 5627 17370 5727
rect 16919 5275 17019 5627
rect 13848 5175 17019 5275
rect 17711 5175 20595 5275
rect 13848 4659 14261 4759
rect 14161 3717 14261 4659
rect 11817 3617 14261 3717
rect 11817 195 11917 3617
rect 15679 195 15779 5175
rect 17711 5081 17811 5175
rect 17373 4981 17811 5081
rect 19548 195 19648 5175
rect 20245 4659 20595 4759
rect 20245 3723 20345 4659
rect 20245 3623 23511 3723
rect 23411 195 23511 3623
rect 27274 195 27374 8277
rect 7910 25 7919 195
rect 8089 25 8098 195
rect 11774 25 11783 195
rect 11953 25 11962 195
rect 15638 25 15647 195
rect 15817 25 15826 195
rect 19502 25 19511 195
rect 19681 25 19690 195
rect 23366 25 23375 195
rect 23545 25 23554 195
rect 27230 25 27239 195
rect 27409 25 27418 195
<< via2 >>
rect 3006 44614 3066 44674
rect 3558 44614 3618 44674
rect 4110 44614 4170 44674
rect 4662 44614 4722 44674
rect 5214 44614 5274 44674
rect 5766 44614 5826 44674
rect 6318 44614 6378 44674
rect 6870 44614 6930 44674
rect 7422 44614 7482 44674
rect 7974 44614 8034 44674
rect 8526 44614 8586 44674
rect 9078 44614 9138 44674
rect 9630 44614 9690 44674
rect 10182 44614 10242 44674
rect 10734 44614 10794 44674
rect 11286 44614 11346 44674
rect 11838 44614 11898 44674
rect 12390 44614 12450 44674
rect 12942 44614 13002 44674
rect 13494 44614 13554 44674
rect 14046 44614 14106 44674
rect 14598 44614 14658 44674
rect 15150 44614 15210 44674
rect 15702 44614 15762 44674
rect 20670 44614 20730 44674
rect 21222 44614 21282 44674
rect 21774 44614 21834 44674
rect 22326 44614 22386 44674
rect 22878 44614 22938 44674
rect 23430 44614 23490 44674
rect 23982 44614 24042 44674
rect 24534 44614 24594 44674
rect 7919 25 8089 195
rect 11783 25 11953 195
rect 15647 25 15817 195
rect 19511 25 19681 195
rect 23375 25 23545 195
rect 27239 25 27409 195
<< metal3 >>
rect 3001 45016 3071 45017
rect 3553 45016 3623 45017
rect 4105 45016 4175 45017
rect 4657 45016 4727 45017
rect 5209 45016 5279 45017
rect 5761 45016 5831 45017
rect 6313 45016 6383 45017
rect 6865 45016 6935 45017
rect 7417 45016 7487 45017
rect 7969 45016 8039 45017
rect 8521 45016 8591 45017
rect 9073 45016 9143 45017
rect 9625 45016 9695 45017
rect 10177 45016 10247 45017
rect 10729 45016 10799 45017
rect 11281 45016 11351 45017
rect 11833 45016 11903 45017
rect 12385 45016 12455 45017
rect 12937 45016 13007 45017
rect 13489 45016 13559 45017
rect 14041 45016 14111 45017
rect 14593 45016 14663 45017
rect 15145 45016 15215 45017
rect 15697 45016 15767 45017
rect 20665 45016 20735 45017
rect 21217 45016 21287 45017
rect 21769 45016 21839 45017
rect 22321 45016 22391 45017
rect 22873 45016 22943 45017
rect 23425 45016 23495 45017
rect 23977 45016 24047 45017
rect 24529 45016 24599 45017
rect 2996 44948 3002 45016
rect 3070 44948 3076 45016
rect 3548 44948 3554 45016
rect 3622 44948 3628 45016
rect 4100 44948 4106 45016
rect 4174 44948 4180 45016
rect 4652 44948 4658 45016
rect 4726 44948 4732 45016
rect 5204 44948 5210 45016
rect 5278 44948 5284 45016
rect 5756 44948 5762 45016
rect 5830 44948 5836 45016
rect 6308 44948 6314 45016
rect 6382 44948 6388 45016
rect 6860 44948 6866 45016
rect 6934 44948 6940 45016
rect 7412 44948 7418 45016
rect 7486 44948 7492 45016
rect 7964 44948 7970 45016
rect 8038 44948 8044 45016
rect 8516 44948 8522 45016
rect 8590 44948 8596 45016
rect 9068 44948 9074 45016
rect 9142 44948 9148 45016
rect 9620 44948 9626 45016
rect 9694 44948 9700 45016
rect 10172 44948 10178 45016
rect 10246 44948 10252 45016
rect 10724 44948 10730 45016
rect 10798 44948 10804 45016
rect 11276 44948 11282 45016
rect 11350 44948 11356 45016
rect 11828 44948 11834 45016
rect 11902 44948 11908 45016
rect 12380 44948 12386 45016
rect 12454 44948 12460 45016
rect 12932 44948 12938 45016
rect 13006 44948 13012 45016
rect 13484 44948 13490 45016
rect 13558 44948 13564 45016
rect 14036 44948 14042 45016
rect 14110 44948 14116 45016
rect 14588 44948 14594 45016
rect 14662 44948 14668 45016
rect 15140 44948 15146 45016
rect 15214 44948 15220 45016
rect 15692 44948 15698 45016
rect 15766 44948 15772 45016
rect 20660 44948 20666 45016
rect 20734 44948 20740 45016
rect 21212 44948 21218 45016
rect 21286 44948 21292 45016
rect 21764 44948 21770 45016
rect 21838 44948 21844 45016
rect 22316 44948 22322 45016
rect 22390 44948 22396 45016
rect 22868 44948 22874 45016
rect 22942 44948 22948 45016
rect 23420 44948 23426 45016
rect 23494 44948 23500 45016
rect 23972 44948 23978 45016
rect 24046 44948 24052 45016
rect 24524 44948 24530 45016
rect 24598 44948 24604 45016
rect 3001 44674 3071 44948
rect 3001 44614 3006 44674
rect 3066 44614 3071 44674
rect 3001 44607 3071 44614
rect 3553 44674 3623 44948
rect 3553 44614 3558 44674
rect 3618 44614 3623 44674
rect 3553 44607 3623 44614
rect 4105 44674 4175 44948
rect 4105 44614 4110 44674
rect 4170 44614 4175 44674
rect 4105 44607 4175 44614
rect 4657 44674 4727 44948
rect 4657 44614 4662 44674
rect 4722 44614 4727 44674
rect 4657 44607 4727 44614
rect 5209 44674 5279 44948
rect 5209 44614 5214 44674
rect 5274 44614 5279 44674
rect 5209 44607 5279 44614
rect 5761 44674 5831 44948
rect 5761 44614 5766 44674
rect 5826 44614 5831 44674
rect 5761 44607 5831 44614
rect 6313 44674 6383 44948
rect 6313 44614 6318 44674
rect 6378 44614 6383 44674
rect 6313 44607 6383 44614
rect 6865 44674 6935 44948
rect 6865 44614 6870 44674
rect 6930 44614 6935 44674
rect 6865 44607 6935 44614
rect 7417 44674 7487 44948
rect 7417 44614 7422 44674
rect 7482 44614 7487 44674
rect 7417 44607 7487 44614
rect 7969 44674 8039 44948
rect 7969 44614 7974 44674
rect 8034 44614 8039 44674
rect 7969 44607 8039 44614
rect 8521 44674 8591 44948
rect 8521 44614 8526 44674
rect 8586 44614 8591 44674
rect 8521 44607 8591 44614
rect 9073 44674 9143 44948
rect 9073 44614 9078 44674
rect 9138 44614 9143 44674
rect 9073 44607 9143 44614
rect 9625 44674 9695 44948
rect 9625 44614 9630 44674
rect 9690 44614 9695 44674
rect 9625 44607 9695 44614
rect 10177 44674 10247 44948
rect 10177 44614 10182 44674
rect 10242 44614 10247 44674
rect 10177 44607 10247 44614
rect 10729 44674 10799 44948
rect 10729 44614 10734 44674
rect 10794 44614 10799 44674
rect 10729 44607 10799 44614
rect 11281 44674 11351 44948
rect 11281 44614 11286 44674
rect 11346 44614 11351 44674
rect 11281 44607 11351 44614
rect 11833 44674 11903 44948
rect 11833 44614 11838 44674
rect 11898 44614 11903 44674
rect 11833 44607 11903 44614
rect 12385 44674 12455 44948
rect 12385 44614 12390 44674
rect 12450 44614 12455 44674
rect 12385 44607 12455 44614
rect 12937 44674 13007 44948
rect 12937 44614 12942 44674
rect 13002 44614 13007 44674
rect 12937 44607 13007 44614
rect 13489 44674 13559 44948
rect 13489 44614 13494 44674
rect 13554 44614 13559 44674
rect 13489 44607 13559 44614
rect 14041 44674 14111 44948
rect 14041 44614 14046 44674
rect 14106 44614 14111 44674
rect 14041 44607 14111 44614
rect 14593 44674 14663 44948
rect 14593 44614 14598 44674
rect 14658 44614 14663 44674
rect 14593 44607 14663 44614
rect 15145 44674 15215 44948
rect 15145 44614 15150 44674
rect 15210 44614 15215 44674
rect 15145 44607 15215 44614
rect 15697 44674 15767 44948
rect 15697 44614 15702 44674
rect 15762 44614 15767 44674
rect 15697 44607 15767 44614
rect 20665 44674 20735 44948
rect 20665 44614 20670 44674
rect 20730 44614 20735 44674
rect 20665 44607 20735 44614
rect 21217 44674 21287 44948
rect 21217 44614 21222 44674
rect 21282 44614 21287 44674
rect 21217 44607 21287 44614
rect 21769 44674 21839 44948
rect 21769 44614 21774 44674
rect 21834 44614 21839 44674
rect 21769 44607 21839 44614
rect 22321 44674 22391 44948
rect 22321 44614 22326 44674
rect 22386 44614 22391 44674
rect 22321 44607 22391 44614
rect 22873 44674 22943 44948
rect 22873 44614 22878 44674
rect 22938 44614 22943 44674
rect 22873 44607 22943 44614
rect 23425 44674 23495 44948
rect 23425 44614 23430 44674
rect 23490 44614 23495 44674
rect 23425 44607 23495 44614
rect 23977 44674 24047 44948
rect 23977 44614 23982 44674
rect 24042 44614 24047 44674
rect 23977 44607 24047 44614
rect 24529 44674 24599 44948
rect 24529 44614 24534 44674
rect 24594 44614 24599 44674
rect 24529 44607 24599 44614
rect 7914 199 8094 200
rect 11778 199 11958 200
rect 15642 199 15822 200
rect 19506 199 19686 200
rect 23370 199 23550 200
rect 27234 199 27414 200
rect 7909 21 7915 199
rect 8093 21 8099 199
rect 11773 21 11779 199
rect 11957 21 11963 199
rect 15637 21 15643 199
rect 15821 21 15827 199
rect 19501 21 19507 199
rect 19685 21 19691 199
rect 23365 21 23371 199
rect 23549 21 23555 199
rect 27229 21 27235 199
rect 27413 21 27419 199
rect 7914 20 8094 21
rect 11778 20 11958 21
rect 15642 20 15822 21
rect 19506 20 19686 21
rect 23370 20 23550 21
rect 27234 20 27414 21
<< via3 >>
rect 3002 44948 3070 45016
rect 3554 44948 3622 45016
rect 4106 44948 4174 45016
rect 4658 44948 4726 45016
rect 5210 44948 5278 45016
rect 5762 44948 5830 45016
rect 6314 44948 6382 45016
rect 6866 44948 6934 45016
rect 7418 44948 7486 45016
rect 7970 44948 8038 45016
rect 8522 44948 8590 45016
rect 9074 44948 9142 45016
rect 9626 44948 9694 45016
rect 10178 44948 10246 45016
rect 10730 44948 10798 45016
rect 11282 44948 11350 45016
rect 11834 44948 11902 45016
rect 12386 44948 12454 45016
rect 12938 44948 13006 45016
rect 13490 44948 13558 45016
rect 14042 44948 14110 45016
rect 14594 44948 14662 45016
rect 15146 44948 15214 45016
rect 15698 44948 15766 45016
rect 20666 44948 20734 45016
rect 21218 44948 21286 45016
rect 21770 44948 21838 45016
rect 22322 44948 22390 45016
rect 22874 44948 22942 45016
rect 23426 44948 23494 45016
rect 23978 44948 24046 45016
rect 24530 44948 24598 45016
rect 7915 195 8093 199
rect 7915 25 7919 195
rect 7919 25 8089 195
rect 8089 25 8093 195
rect 7915 21 8093 25
rect 11779 195 11957 199
rect 11779 25 11783 195
rect 11783 25 11953 195
rect 11953 25 11957 195
rect 11779 21 11957 25
rect 15643 195 15821 199
rect 15643 25 15647 195
rect 15647 25 15817 195
rect 15817 25 15821 195
rect 15643 21 15821 25
rect 19507 195 19685 199
rect 19507 25 19511 195
rect 19511 25 19681 195
rect 19681 25 19685 195
rect 19507 21 19685 25
rect 23371 195 23549 199
rect 23371 25 23375 195
rect 23375 25 23545 195
rect 23545 25 23549 195
rect 23371 21 23549 25
rect 27235 195 27413 199
rect 27235 25 27239 195
rect 27239 25 27409 195
rect 27409 25 27413 195
rect 27235 21 27413 25
<< metal4 >>
rect 3006 45017 3066 45152
rect 3558 45017 3618 45152
rect 4110 45018 4170 45152
rect 4107 45017 4173 45018
rect 4662 45017 4722 45152
rect 5214 45017 5274 45152
rect 5766 45017 5826 45152
rect 6318 45017 6378 45152
rect 6870 45017 6930 45152
rect 7422 45017 7482 45152
rect 7974 45017 8034 45152
rect 8526 45017 8586 45152
rect 9078 45017 9138 45152
rect 9630 45017 9690 45152
rect 10182 45017 10242 45152
rect 10734 45017 10794 45152
rect 11286 45017 11346 45152
rect 11838 45017 11898 45152
rect 12390 45017 12450 45152
rect 12942 45017 13002 45152
rect 13494 45017 13554 45152
rect 14046 45017 14106 45152
rect 14598 45017 14658 45152
rect 15150 45017 15210 45152
rect 15702 45017 15762 45152
rect 3001 45016 3071 45017
rect 3001 44948 3002 45016
rect 3070 44948 3071 45016
rect 3001 44947 3071 44948
rect 3553 45016 3623 45017
rect 3553 44948 3554 45016
rect 3622 44948 3623 45016
rect 3553 44947 3623 44948
rect 4105 45016 4175 45017
rect 4105 44948 4106 45016
rect 4174 44948 4175 45016
rect 4105 44947 4175 44948
rect 4657 45016 4727 45017
rect 4657 44948 4658 45016
rect 4726 44948 4727 45016
rect 4657 44947 4727 44948
rect 5209 45016 5279 45017
rect 5209 44948 5210 45016
rect 5278 44948 5279 45016
rect 5209 44947 5279 44948
rect 5761 45016 5831 45017
rect 5761 44948 5762 45016
rect 5830 44948 5831 45016
rect 5761 44947 5831 44948
rect 6313 45016 6383 45017
rect 6313 44948 6314 45016
rect 6382 44948 6383 45016
rect 6313 44947 6383 44948
rect 6865 45016 6935 45017
rect 6865 44948 6866 45016
rect 6934 44948 6935 45016
rect 6865 44947 6935 44948
rect 7417 45016 7487 45017
rect 7417 44948 7418 45016
rect 7486 44948 7487 45016
rect 7417 44947 7487 44948
rect 7969 45016 8039 45017
rect 7969 44948 7970 45016
rect 8038 44948 8039 45016
rect 7969 44947 8039 44948
rect 8521 45016 8591 45017
rect 8521 44948 8522 45016
rect 8590 44948 8591 45016
rect 8521 44947 8591 44948
rect 9073 45016 9143 45017
rect 9073 44948 9074 45016
rect 9142 44948 9143 45016
rect 9073 44947 9143 44948
rect 9625 45016 9695 45017
rect 9625 44948 9626 45016
rect 9694 44948 9695 45016
rect 9625 44947 9695 44948
rect 10177 45016 10247 45017
rect 10177 44948 10178 45016
rect 10246 44948 10247 45016
rect 10177 44947 10247 44948
rect 10729 45016 10799 45017
rect 10729 44948 10730 45016
rect 10798 44948 10799 45016
rect 10729 44947 10799 44948
rect 11281 45016 11351 45017
rect 11281 44948 11282 45016
rect 11350 44948 11351 45016
rect 11281 44947 11351 44948
rect 11833 45016 11903 45017
rect 11833 44948 11834 45016
rect 11902 44948 11903 45016
rect 11833 44947 11903 44948
rect 12385 45016 12455 45017
rect 12385 44948 12386 45016
rect 12454 44948 12455 45016
rect 12385 44947 12455 44948
rect 12937 45016 13007 45017
rect 12937 44948 12938 45016
rect 13006 44948 13007 45016
rect 12937 44947 13007 44948
rect 13489 45016 13559 45017
rect 13489 44948 13490 45016
rect 13558 44948 13559 45016
rect 13489 44947 13559 44948
rect 14041 45016 14111 45017
rect 14041 44948 14042 45016
rect 14110 44948 14111 45016
rect 14041 44947 14111 44948
rect 14593 45016 14663 45017
rect 14593 44948 14594 45016
rect 14662 44948 14663 45016
rect 14593 44947 14663 44948
rect 15145 45016 15215 45017
rect 15145 44948 15146 45016
rect 15214 44948 15215 45016
rect 15145 44947 15215 44948
rect 15697 45016 15767 45017
rect 15697 44948 15698 45016
rect 15766 44948 15767 45016
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 45017 19626 45152
rect 19566 44952 19631 45017
rect 20118 44952 20178 45152
rect 20670 45017 20730 45152
rect 21222 45017 21282 45152
rect 21774 45017 21834 45152
rect 22326 45017 22386 45152
rect 22878 45017 22938 45152
rect 23430 45017 23490 45152
rect 23982 45017 24042 45152
rect 24534 45017 24594 45152
rect 20665 45016 20735 45017
rect 15697 44947 15767 44948
rect 20665 44948 20666 45016
rect 20734 44948 20735 45016
rect 20665 44947 20735 44948
rect 21217 45016 21287 45017
rect 21217 44948 21218 45016
rect 21286 44948 21287 45016
rect 21217 44947 21287 44948
rect 21769 45016 21839 45017
rect 21769 44948 21770 45016
rect 21838 44948 21839 45016
rect 21769 44947 21839 44948
rect 22321 45016 22391 45017
rect 22321 44948 22322 45016
rect 22390 44948 22391 45016
rect 22321 44947 22391 44948
rect 22873 45016 22943 45017
rect 22873 44948 22874 45016
rect 22942 44948 22943 45016
rect 22873 44947 22943 44948
rect 23425 45016 23495 45017
rect 23425 44948 23426 45016
rect 23494 44948 23495 45016
rect 23425 44947 23495 44948
rect 23977 45016 24047 45017
rect 23977 44948 23978 45016
rect 24046 44948 24047 45016
rect 23977 44947 24047 44948
rect 24529 45016 24599 45017
rect 24529 44948 24530 45016
rect 24598 44948 24599 45016
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 24529 44947 24599 44948
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 199 8094 200
rect 7914 21 7915 199
rect 8093 21 8094 199
rect 7914 0 8094 21
rect 11778 199 11958 200
rect 11778 21 11779 199
rect 11957 21 11958 199
rect 11778 0 11958 21
rect 15642 199 15822 200
rect 15642 21 15643 199
rect 15821 21 15822 199
rect 15642 0 15822 21
rect 19506 199 19686 200
rect 19506 21 19507 199
rect 19685 21 19686 199
rect 19506 0 19686 21
rect 23370 199 23550 200
rect 23370 21 23371 199
rect 23549 21 23550 199
rect 23370 0 23550 21
rect 27234 199 27414 200
rect 27234 21 27235 199
rect 27413 21 27414 199
rect 27234 0 27414 21
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
