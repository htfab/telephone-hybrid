magic
tech sky130A
magscale 1 2
timestamp 1731102314
<< dnwell >>
rect -438 -275 4076 10803
<< nwell >>
rect -518 10597 4156 10883
rect -518 -69 -232 10597
rect 3870 -69 4156 10597
rect -518 -355 4156 -69
<< nsubdiff >>
rect -481 10826 4119 10846
rect -481 10792 -401 10826
rect 4039 10792 4119 10826
rect -481 10772 4119 10792
rect -481 10766 -407 10772
rect -481 -238 -461 10766
rect -427 -238 -407 10766
rect -481 -244 -407 -238
rect 4045 10766 4119 10772
rect 4045 -238 4065 10766
rect 4099 -238 4119 10766
rect 4045 -244 4119 -238
rect -481 -264 4119 -244
rect -481 -298 -401 -264
rect 4039 -298 4119 -264
rect -481 -318 4119 -298
<< nsubdiffcont >>
rect -401 10792 4039 10826
rect -461 -238 -427 10766
rect 4065 -238 4099 10766
rect -401 -298 4039 -264
<< locali >>
rect -461 10792 -401 10826
rect 4039 10792 4099 10826
rect -461 10766 -427 10792
rect -461 -264 -427 -238
rect 4065 10766 4099 10792
rect 4065 -264 4099 -238
rect -461 -298 -401 -264
rect 4039 -298 4099 -264
use hybrid  hybrid_0
timestamp 1727597281
transform 1 0 -3204 0 1 3276
box 3204 -3276 7092 7391
<< end >>
