magic
tech sky130A
magscale 1 2
timestamp 1727637087
<< nwell >>
rect -60 606 2636 1292
<< pwell >>
rect -60 556 126 557
rect -60 0 2636 556
<< mvpsubdiff >>
rect -14 508 2600 520
rect -14 474 124 508
rect 352 474 424 508
rect 652 474 724 508
rect 952 474 1024 508
rect 1252 474 1324 508
rect 1552 474 1624 508
rect 1852 474 1924 508
rect 2152 474 2224 508
rect 2452 474 2600 508
rect -14 462 2600 474
rect -14 412 44 462
rect -14 144 -2 412
rect 32 144 44 412
rect -14 94 44 144
rect 2542 412 2600 462
rect 2542 144 2554 412
rect 2588 144 2600 412
rect 2542 94 2600 144
rect -14 82 2600 94
rect -14 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2600 82
rect -14 36 2600 48
<< mvnsubdiff >>
rect 6 1214 2570 1226
rect 6 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2570 1214
rect 6 1168 2570 1180
rect 6 1118 64 1168
rect 6 780 18 1118
rect 52 780 64 1118
rect 6 730 64 780
rect 2512 1118 2570 1168
rect 2512 780 2524 1118
rect 2558 780 2570 1118
rect 2512 730 2570 780
rect 6 718 2570 730
rect 6 684 124 718
rect 352 684 424 718
rect 652 684 724 718
rect 952 684 1024 718
rect 1252 684 1324 718
rect 1552 684 1624 718
rect 1852 684 1924 718
rect 2152 684 2224 718
rect 2452 684 2570 718
rect 6 672 2570 684
<< mvpsubdiffcont >>
rect 124 474 352 508
rect 424 474 652 508
rect 724 474 952 508
rect 1024 474 1252 508
rect 1324 474 1552 508
rect 1624 474 1852 508
rect 1924 474 2152 508
rect 2224 474 2452 508
rect -2 144 32 412
rect 2554 144 2588 412
rect 124 48 352 82
rect 424 48 652 82
rect 724 48 952 82
rect 1024 48 1252 82
rect 1324 48 1552 82
rect 1624 48 1852 82
rect 1924 48 2152 82
rect 2224 48 2452 82
<< mvnsubdiffcont >>
rect 124 1180 352 1214
rect 424 1180 652 1214
rect 724 1180 952 1214
rect 1024 1180 1252 1214
rect 1324 1180 1552 1214
rect 1624 1180 1852 1214
rect 1924 1180 2152 1214
rect 2224 1180 2452 1214
rect 18 780 52 1118
rect 2524 780 2558 1118
rect 124 684 352 718
rect 424 684 652 718
rect 724 684 952 718
rect 1024 684 1252 718
rect 1324 684 1552 718
rect 1624 684 1852 718
rect 1924 684 2152 718
rect 2224 684 2452 718
<< locali >>
rect 18 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2558 1214
rect 18 1118 52 1180
rect 18 718 52 780
rect 2524 1118 2558 1180
rect 2524 718 2558 780
rect 18 684 124 718
rect 352 684 424 718
rect 652 684 724 718
rect 952 684 1024 718
rect 1252 684 1324 718
rect 1552 684 1624 718
rect 1852 684 1924 718
rect 2152 684 2224 718
rect 2452 684 2558 718
rect -2 474 124 508
rect 352 474 424 508
rect 652 474 724 508
rect 952 474 1024 508
rect 1252 474 1324 508
rect 1552 474 1624 508
rect 1852 474 1924 508
rect 2152 474 2224 508
rect 2452 474 2588 508
rect -2 412 32 474
rect -2 82 32 144
rect 2554 412 2588 474
rect 2554 82 2588 144
rect -2 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2588 82
<< viali >>
rect 124 1180 352 1214
rect 424 1180 652 1214
rect 724 1180 952 1214
rect 1024 1180 1252 1214
rect 1324 1180 1552 1214
rect 1624 1180 1852 1214
rect 1924 1180 2152 1214
rect 2224 1180 2452 1214
rect 124 48 352 82
rect 424 48 652 82
rect 724 48 952 82
rect 1024 48 1252 82
rect 1324 48 1552 82
rect 1624 48 1852 82
rect 1924 48 2152 82
rect 2224 48 2452 82
<< metal1 >>
rect 88 1214 2488 1226
rect 88 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2488 1214
rect 88 1168 2488 1180
rect 88 82 2488 94
rect 88 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2488 82
rect 88 36 2488 48
<< labels >>
flabel metal1 88 1168 2488 1226 0 FreeSans 256 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal1 88 36 2488 94 0 FreeSans 256 0 0 0 VSS
port 1 nsew ground bidirectional
<< end >>
