magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< nwell >>
rect 0 954 476 2076
<< pwell >>
rect 0 0 476 904
<< mvpsubdiff >>
rect 100 856 376 868
rect 100 822 124 856
rect 352 822 376 856
rect 100 810 376 822
rect 100 82 376 94
rect 100 48 124 82
rect 352 48 376 82
rect 100 36 376 48
<< mvnsubdiff >>
rect 100 1998 376 2010
rect 100 1964 124 1998
rect 352 1964 376 1998
rect 100 1952 376 1964
rect 100 1066 376 1078
rect 100 1032 124 1066
rect 352 1032 376 1066
rect 100 1020 376 1032
<< mvpsubdiffcont >>
rect 124 822 352 856
rect 124 48 352 82
<< mvnsubdiffcont >>
rect 124 1964 352 1998
rect 124 1032 352 1066
<< locali >>
rect 100 1964 124 1998
rect 352 1964 376 1998
rect 100 1032 124 1066
rect 352 1032 376 1066
rect 100 822 124 856
rect 352 822 376 856
rect 100 48 124 82
rect 352 48 376 82
<< viali >>
rect 204 1964 272 1998
rect 204 48 272 82
<< metal1 >>
rect 118 1952 124 2004
rect 250 1998 284 2004
rect 272 1964 284 1998
rect 250 1958 284 1964
rect 250 1952 256 1958
rect 118 1633 164 1952
rect 215 1595 261 1900
rect 192 1543 204 1595
rect 272 1543 284 1595
rect 112 1492 164 1498
rect 312 1484 358 1834
rect 112 1434 164 1440
rect 118 679 164 1434
rect 215 1165 261 1464
rect 272 1438 358 1484
rect 312 1326 358 1398
rect 352 1220 358 1326
rect 300 1209 358 1220
rect 192 1159 284 1165
rect 192 1107 204 1159
rect 272 1107 284 1159
rect 192 1101 284 1107
rect 192 720 204 772
rect 272 720 284 772
rect 118 573 124 679
rect 118 561 164 573
rect 215 505 261 720
rect 312 561 358 1209
rect 250 399 261 505
rect 118 94 164 343
rect 215 155 261 399
rect 312 331 358 343
rect 352 225 358 331
rect 312 213 358 225
rect 118 42 124 94
rect 250 88 256 94
rect 250 82 284 88
rect 272 48 284 82
rect 250 42 284 48
<< via1 >>
rect 124 1998 250 2004
rect 124 1964 204 1998
rect 204 1964 250 1998
rect 124 1952 250 1964
rect 204 1543 272 1595
rect 112 1440 164 1492
rect 300 1220 352 1326
rect 204 1107 272 1159
rect 204 720 272 772
rect 124 573 176 679
rect 198 399 250 505
rect 300 225 352 331
rect 124 82 250 94
rect 124 48 204 82
rect 204 48 250 82
rect 124 42 250 48
<< metal2 >>
rect 118 1952 124 2004
rect 250 1952 256 2004
rect 118 1866 256 1952
rect 118 1649 256 1787
rect 118 1498 164 1649
rect 192 1595 358 1601
rect 192 1543 204 1595
rect 272 1543 358 1595
rect 192 1537 358 1543
rect 112 1492 164 1498
rect 112 1434 164 1440
rect 215 1463 358 1537
rect 215 1406 261 1463
rect 118 1360 261 1406
rect 118 769 164 1360
rect 220 1326 358 1332
rect 220 1220 300 1326
rect 352 1220 358 1326
rect 220 1193 358 1220
rect 192 1159 284 1165
rect 192 1107 204 1159
rect 272 1156 284 1159
rect 272 1110 358 1156
rect 272 1107 284 1110
rect 192 1101 284 1107
rect 192 772 284 778
rect 192 769 204 772
rect 118 723 204 769
rect 192 720 204 723
rect 272 720 284 772
rect 192 714 284 720
rect 118 679 256 685
rect 118 573 124 679
rect 176 573 256 679
rect 118 547 256 573
rect 118 505 256 513
rect 118 399 198 505
rect 250 399 256 505
rect 118 375 256 399
rect 312 343 358 1110
rect 294 331 358 343
rect 294 225 300 331
rect 352 225 358 331
rect 294 213 358 225
rect 118 94 256 180
rect 118 42 124 94
rect 250 42 256 94
use sky130_fd_pr__nfet_g5v0d10v5_83EA8U  sky130_fd_pr__nfet_g5v0d10v5_83EA8U_0
timestamp 1727597281
transform 1 0 238 0 1 452
box -108 -327 108 327
use sky130_fd_pr__pfet_g5v0d10v5_KLSDQ5  sky130_fd_pr__pfet_g5v0d10v5_KLSDQ5_1
timestamp 1727597281
transform 1 0 238 0 1 1515
box -174 -418 174 418
<< labels >>
flabel metal2 118 375 256 513 0 FreeSans 256 0 0 0 EN
port 0 nsew
flabel metal2 118 547 256 685 0 FreeSans 256 0 0 0 UA
port 1 nsew
flabel metal2 220 1193 358 1331 0 FreeSans 256 0 0 0 UB
port 2 nsew
flabel metal2 118 1866 256 2004 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal2 118 42 256 180 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
