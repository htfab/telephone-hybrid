magic
tech sky130A
magscale 1 2
timestamp 1731100676
<< metal1 >>
rect 3074 11099 3212 11105
rect 3212 10961 7414 11099
rect 3074 10955 3212 10961
rect 3074 9887 3212 9893
rect 3212 9749 7414 9887
rect 3074 9743 3212 9749
rect 3074 1705 3212 1711
rect 3212 1567 7414 1705
rect 3074 1561 3212 1567
rect 3074 493 3212 499
rect 3212 355 7414 493
rect 3074 349 3212 355
<< via1 >>
rect 3074 10961 3212 11099
rect 3074 9749 3212 9887
rect 3074 1567 3212 1705
rect 3074 355 3212 493
<< metal2 >>
rect 4644 11874 4678 12445
rect 4504 11840 4678 11874
rect 4365 11622 4425 11631
rect 4504 11609 4538 11840
rect 4425 11575 4538 11609
rect 4630 11714 4690 11748
rect 4365 11553 4425 11562
rect 4239 11496 4299 11505
rect 4630 11483 4664 11714
rect 4299 11449 4664 11483
rect 4239 11427 4299 11436
rect 277 11273 415 11411
rect 2761 11273 3212 11411
rect 3074 11099 3212 11273
rect 4617 11116 4677 11125
rect 3068 10961 3074 11099
rect 3212 10961 3218 11099
rect 4617 11047 4677 11056
rect 4491 10419 4551 10428
rect 4551 10372 4678 10406
rect 4491 10350 4551 10359
rect 4113 10293 4173 10302
rect 4617 10293 4677 10302
rect 4173 10246 4617 10280
rect 4113 10224 4173 10233
rect 4617 10224 4677 10233
rect 3987 10167 4047 10176
rect 4491 10167 4551 10176
rect 4047 10120 4491 10154
rect 3987 10098 4047 10107
rect 4491 10098 4551 10107
rect 3068 9749 3074 9887
rect 3212 9749 3218 9887
rect 4617 9774 4677 9783
rect 3074 9587 3212 9749
rect 4617 9705 4677 9714
rect 2761 9449 3212 9587
rect 4491 9077 4551 9086
rect 4551 9030 4678 9064
rect 4491 9008 4551 9017
rect 4365 8432 4425 8441
rect 4425 8385 4678 8419
rect 4365 8363 4425 8372
rect 4239 7735 4299 7744
rect 4299 7688 4678 7722
rect 4239 7666 4299 7675
rect 3735 7090 3795 7099
rect 3795 7043 4678 7077
rect 3735 7021 3795 7030
rect 3861 6393 3921 6402
rect 3921 6346 4678 6380
rect 3861 6324 3921 6333
rect 4617 5748 4677 5757
rect 4617 5679 4677 5688
rect 4491 5051 4551 5060
rect 4551 5004 4678 5038
rect 4491 4982 4551 4991
rect 4239 4406 4299 4415
rect 4299 4359 4678 4393
rect 4239 4337 4299 4346
rect 4365 3709 4425 3718
rect 4425 3662 4678 3696
rect 6990 3662 7867 3696
rect 4365 3640 4425 3649
rect 3987 3064 4047 3073
rect 4047 3017 4678 3051
rect 3987 2995 4047 3004
rect 4113 2367 4173 2376
rect 4173 2320 4678 2354
rect 6990 2320 7867 2354
rect 4113 2298 4173 2307
rect 2760 1866 3212 2004
rect 3074 1705 3212 1866
rect 3068 1567 3074 1705
rect 3212 1567 3218 1705
rect 6990 978 7867 1012
rect 3068 355 3074 493
rect 3212 355 3218 493
rect 3074 180 3212 355
rect 276 42 414 180
rect 2760 42 3212 180
rect 6990 -364 7867 -330
<< via2 >>
rect 4365 11562 4425 11622
rect 4239 11436 4299 11496
rect 4617 11056 4677 11116
rect 4491 10359 4551 10419
rect 4113 10233 4173 10293
rect 4617 10233 4677 10293
rect 3987 10107 4047 10167
rect 4491 10107 4551 10167
rect 4617 9714 4677 9774
rect 4491 9017 4551 9077
rect 4365 8372 4425 8432
rect 4239 7675 4299 7735
rect 3735 7030 3795 7090
rect 3861 6333 3921 6393
rect 4617 5688 4677 5748
rect 4491 4991 4551 5051
rect 4239 4346 4299 4406
rect 4365 3649 4425 3709
rect 3987 3004 4047 3064
rect 4113 2307 4173 2367
rect 562 569 680 679
<< metal3 >>
rect 694 11814 4677 11874
rect 694 10909 754 11814
rect 970 11688 4551 11748
rect 970 10909 1030 11688
rect 4360 11622 4430 11627
rect 1246 11562 4365 11622
rect 4425 11562 4430 11622
rect 1246 10909 1306 11562
rect 4360 11557 4430 11562
rect 4234 11496 4304 11501
rect 1522 11436 4239 11496
rect 4299 11436 4304 11496
rect 1522 10909 1582 11436
rect 4234 11431 4304 11436
rect 1798 11310 4425 11370
rect 1798 10909 1858 11310
rect 2074 11184 4299 11244
rect 2074 10909 2134 11184
rect 2350 11058 4173 11118
rect 2350 10909 2410 11058
rect 2626 10909 4047 10969
rect 3987 10172 4047 10909
rect 4113 10298 4173 11058
rect 4108 10293 4178 10298
rect 4108 10233 4113 10293
rect 4173 10233 4178 10293
rect 4108 10228 4178 10233
rect 3982 10167 4052 10172
rect 3982 10107 3987 10167
rect 4047 10107 4052 10167
rect 3982 10102 4052 10107
rect 4239 7740 4299 11184
rect 4365 8437 4425 11310
rect 4491 10424 4551 11688
rect 4617 11121 4677 11814
rect 4612 11116 4682 11121
rect 4612 11056 4617 11116
rect 4677 11056 4682 11116
rect 4612 11051 4682 11056
rect 4486 10419 4556 10424
rect 4486 10359 4491 10419
rect 4551 10359 4556 10419
rect 4486 10354 4556 10359
rect 4612 10293 4682 10298
rect 4612 10233 4617 10293
rect 4677 10233 4682 10293
rect 4612 10228 4682 10233
rect 4486 10167 4556 10172
rect 4486 10107 4491 10167
rect 4551 10107 4556 10167
rect 4486 10102 4556 10107
rect 4491 9082 4551 10102
rect 4617 9779 4677 10228
rect 4612 9774 4682 9779
rect 4612 9714 4617 9774
rect 4677 9714 4682 9774
rect 4612 9709 4682 9714
rect 4486 9077 4556 9082
rect 4486 9017 4491 9077
rect 4551 9017 4556 9077
rect 4486 9012 4556 9017
rect 4360 8432 4430 8437
rect 4360 8372 4365 8432
rect 4425 8372 4430 8432
rect 4360 8367 4430 8372
rect 4234 7735 4304 7740
rect 4234 7675 4239 7735
rect 4299 7675 4304 7735
rect 4234 7670 4304 7675
rect 3730 7090 3800 7095
rect 3730 7030 3735 7090
rect 3795 7030 3800 7090
rect 3730 7025 3800 7030
rect 2760 1649 2898 1787
rect 654 1193 792 1331
rect 3735 1127 3795 7025
rect 3856 6393 3926 6398
rect 3856 6333 3861 6393
rect 3921 6333 3926 6393
rect 3856 6328 3926 6333
rect 1143 1067 3795 1127
rect 552 679 690 701
rect 552 569 562 679
rect 680 569 690 679
rect 552 563 690 569
rect 591 199 651 474
rect 867 325 927 474
rect 1143 414 1203 1067
rect 3861 1001 3921 6328
rect 4612 5748 4682 5753
rect 4612 5688 4617 5748
rect 4677 5688 4682 5748
rect 4612 5683 4682 5688
rect 4486 5051 4556 5056
rect 4486 4991 4491 5051
rect 4551 4991 4556 5051
rect 4486 4986 4556 4991
rect 4234 4406 4304 4411
rect 4234 4346 4239 4406
rect 4299 4346 4304 4406
rect 4234 4341 4304 4346
rect 3982 3064 4052 3069
rect 3982 3004 3987 3064
rect 4047 3004 4052 3064
rect 3982 2999 4052 3004
rect 1419 941 3921 1001
rect 1419 414 1479 941
rect 3987 875 4047 2999
rect 4108 2367 4178 2372
rect 4108 2307 4113 2367
rect 4173 2307 4178 2367
rect 4108 2302 4178 2307
rect 1695 815 4047 875
rect 1695 414 1755 815
rect 4113 749 4173 2302
rect 1971 689 4173 749
rect 1971 414 2031 689
rect 4239 623 4299 4341
rect 4360 3709 4430 3714
rect 4360 3649 4365 3709
rect 4425 3649 4430 3709
rect 4360 3644 4430 3649
rect 2247 563 4299 623
rect 2247 414 2307 563
rect 4365 474 4425 3644
rect 2523 414 4425 474
rect 4491 325 4551 4986
rect 867 265 4551 325
rect 4617 199 4677 5683
rect 591 139 4677 199
use decoder4_signed  decoder4_signed_0
timestamp 1731100676
transform -1 0 7562 0 1 -943
box -305 0 2996 13410
use digipot_1hot  x2
timestamp 1727641773
transform 1 0 0 0 1 0
box 110 0 4330 11483
<< labels >>
flabel metal2 276 42 414 180 0 FreeSans 128 0 0 0 VSS
port 7 nsew
flabel metal3 552 563 690 701 0 FreeSans 128 0 0 0 A
port 0 nsew
flabel metal3 2760 1649 2898 1787 0 FreeSans 128 0 0 0 B
port 1 nsew
flabel metal3 654 1193 792 1331 0 FreeSans 128 0 0 0 W
port 8 nsew
flabel metal2 277 11273 415 11411 0 FreeSans 128 0 0 0 VDD
port 6 nsew
flabel metal2 6990 -364 7867 -330 0 FreeSans 128 0 0 0 D3
port 5 nsew
flabel metal2 6990 978 7867 1012 0 FreeSans 128 0 0 0 D0
port 2 nsew
flabel metal2 6990 2320 7867 2354 0 FreeSans 128 0 0 0 D1
port 3 nsew
flabel metal2 6990 3662 7867 3696 0 FreeSans 128 0 0 0 D2
port 4 nsew
<< end >>
