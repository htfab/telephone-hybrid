magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< error_p >>
rect -120 -65 -50 65
rect 50 -65 120 65
<< mvnmos >>
rect -50 -65 50 65
<< mvndiff >>
rect -120 53 -50 65
rect -120 -53 -108 53
rect -74 -53 -50 53
rect -120 -65 -50 -53
rect 50 53 120 65
rect 50 -53 74 53
rect 108 -53 120 53
rect 50 -65 120 -53
<< mvndiffc >>
rect -108 -53 -74 53
rect 74 -53 108 53
<< poly >>
rect -50 137 50 153
rect -50 103 -34 137
rect 34 103 50 137
rect -50 65 50 103
rect -50 -103 50 -65
rect -50 -137 -34 -103
rect 34 -137 50 -103
rect -50 -153 50 -137
<< polycont >>
rect -34 103 34 137
rect -34 -137 34 -103
<< locali >>
rect -50 103 -34 137
rect 34 103 50 137
rect -108 53 -74 69
rect -108 -69 -74 -53
rect 74 53 108 69
rect 74 -69 108 -53
rect -50 -137 -34 -103
rect 34 -137 50 -103
<< viali >>
rect -34 103 34 137
rect -108 -53 -74 53
rect 74 -53 108 53
rect -34 -137 34 -103
<< metal1 >>
rect -46 137 46 143
rect -46 103 -34 137
rect 34 103 46 137
rect -46 97 46 103
rect -114 53 -68 65
rect -114 -53 -108 53
rect -74 -53 -68 53
rect -114 -65 -68 -53
rect 68 53 114 65
rect 68 -53 74 53
rect 108 -53 114 53
rect 68 -65 114 -53
rect -46 -103 46 -97
rect -46 -137 -34 -103
rect 34 -137 46 -103
rect -46 -143 46 -137
<< end >>
