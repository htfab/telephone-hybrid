magic
tech sky130A
magscale 1 2
timestamp 1727638007
<< metal1 >>
rect 88 1168 388 1226
rect 130 845 164 1168
rect 130 94 164 347
rect 221 295 255 1130
rect 312 845 346 1053
rect 312 295 346 347
rect 221 261 346 295
rect 221 141 255 261
rect 312 209 346 261
rect 88 36 388 94
<< labels >>
flabel metal1 88 1168 388 1226 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 88 36 388 94 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 312 845 346 1053 0 FreeSans 256 0 0 0 HI
port 0 nsew
<< end >>
