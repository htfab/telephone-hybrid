magic
tech sky130A
timestamp 1727597281
<< nwell >>
rect 144 303 268 646
<< pwell >>
rect 144 0 268 278
<< mvpsubdiff >>
rect 194 231 250 260
rect 221 206 250 231
rect 221 72 227 206
rect 244 72 250 206
rect 221 47 250 72
rect 194 18 250 47
<< mvnsubdiff >>
rect 194 584 235 613
rect 206 559 235 584
rect 206 390 212 559
rect 229 390 235 559
rect 206 365 235 390
rect 194 336 235 365
<< mvpsubdiffcont >>
rect 227 72 244 206
<< mvnsubdiffcont >>
rect 212 390 229 559
<< locali >>
rect 194 590 229 607
rect 212 559 229 590
rect 212 359 229 390
rect 194 342 229 359
rect 194 237 244 254
rect 227 206 244 237
rect 227 41 244 72
rect 194 24 244 41
<< end >>
