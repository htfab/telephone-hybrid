magic
tech sky130A
magscale 1 2
timestamp 1727641004
<< metal1 >>
rect 118 1952 124 2004
rect 250 1958 284 2004
rect 250 1952 256 1958
rect 118 1633 164 1952
rect 215 1595 261 1900
rect 192 1543 204 1595
rect 272 1543 284 1595
rect 112 1492 164 1498
rect 312 1484 358 1834
rect 112 1434 164 1440
rect 118 685 164 1434
rect 215 1438 358 1484
rect 215 1165 261 1438
rect 312 1332 358 1398
rect 294 1326 358 1332
rect 294 1220 300 1326
rect 352 1220 358 1326
rect 294 1214 358 1220
rect 300 1209 358 1214
rect 192 1159 284 1165
rect 192 1107 204 1159
rect 272 1107 284 1159
rect 192 1101 284 1107
rect 192 720 204 772
rect 272 720 284 772
rect 118 679 182 685
rect 118 573 124 679
rect 176 573 182 679
rect 118 567 182 573
rect 118 561 164 567
rect 215 511 261 720
rect 312 561 358 1209
rect 192 505 261 511
rect 192 399 198 505
rect 250 399 261 505
rect 192 393 261 399
rect 118 94 164 343
rect 215 155 261 393
rect 312 337 358 343
rect 294 331 358 337
rect 294 225 300 331
rect 352 225 358 331
rect 294 219 358 225
rect 312 213 358 219
rect 118 42 124 94
rect 250 88 256 94
rect 250 42 284 88
<< via1 >>
rect 124 1952 250 2004
rect 204 1543 272 1595
rect 112 1440 164 1492
rect 300 1220 352 1326
rect 204 1107 272 1159
rect 204 720 272 772
rect 124 573 176 679
rect 198 399 250 505
rect 300 225 352 331
rect 124 42 250 94
<< metal2 >>
rect 118 1952 124 2004
rect 250 1952 256 2004
rect 118 1866 256 1952
rect 118 1649 256 1787
rect 118 1498 164 1649
rect 192 1595 358 1601
rect 192 1543 204 1595
rect 272 1543 358 1595
rect 192 1537 358 1543
rect 112 1492 164 1498
rect 112 1434 164 1440
rect 215 1463 358 1537
rect 215 1406 261 1463
rect 118 1360 261 1406
rect 118 769 164 1360
rect 220 1326 358 1332
rect 220 1220 300 1326
rect 352 1220 358 1326
rect 220 1193 358 1220
rect 192 1159 284 1165
rect 192 1107 204 1159
rect 272 1156 284 1159
rect 272 1110 358 1156
rect 272 1107 284 1110
rect 192 1101 284 1107
rect 192 772 284 778
rect 192 769 204 772
rect 118 723 204 769
rect 192 720 204 723
rect 272 720 284 772
rect 192 714 284 720
rect 118 679 256 685
rect 118 573 124 679
rect 176 573 256 679
rect 118 547 256 573
rect 118 505 256 513
rect 118 399 198 505
rect 250 399 256 505
rect 118 375 256 399
rect 312 343 358 1110
rect 294 331 358 343
rect 294 225 300 331
rect 352 225 358 331
rect 294 213 358 225
rect 118 94 256 180
rect 118 42 124 94
rect 250 42 256 94
<< labels >>
flabel metal2 118 375 256 513 0 FreeSans 256 0 0 0 EN
port 0 nsew
flabel metal2 118 547 256 685 0 FreeSans 256 0 0 0 UA
port 1 nsew
flabel metal2 220 1193 358 1331 0 FreeSans 256 0 0 0 UB
port 2 nsew
flabel metal2 118 1866 256 2004 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal2 118 42 256 180 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
