MACRO hybrid_dnwell
  CLASS BLOCK ;
  FOREIGN hybrid_dnwell ;
  ORIGIN 2.590 1.775 ;
  SIZE 23.370 BY 56.190 ;
  OBS
      LAYER nwell ;
        RECT -2.590 52.985 20.780 54.415 ;
        RECT -2.590 -0.345 -1.160 52.985 ;
        RECT 2.960 16.000 14.640 16.980 ;
        RECT 2.980 6.220 14.640 16.000 ;
        RECT 19.350 -0.345 20.780 52.985 ;
        RECT -2.590 -1.775 20.780 -0.345 ;
      LAYER li1 ;
        RECT -2.305 53.960 20.495 54.130 ;
        RECT -2.305 -1.320 -2.135 53.960 ;
        RECT 0.000 51.175 0.350 53.335 ;
        RECT 0.830 51.175 1.180 53.335 ;
        RECT 1.660 51.175 2.010 53.335 ;
        RECT 2.490 51.175 2.840 53.335 ;
        RECT 3.320 51.175 3.670 53.335 ;
        RECT 4.150 51.175 4.500 53.335 ;
        RECT 4.980 51.175 5.330 53.335 ;
        RECT 5.810 51.175 6.160 53.335 ;
        RECT 6.640 51.175 6.990 53.335 ;
        RECT 7.470 51.175 7.820 53.335 ;
        RECT 8.300 51.175 8.650 53.335 ;
        RECT 9.130 51.175 9.480 53.335 ;
        RECT 9.960 51.175 10.310 53.335 ;
        RECT 10.790 51.175 11.140 53.335 ;
        RECT 11.620 51.175 11.970 53.335 ;
        RECT 12.450 51.175 12.800 53.335 ;
        RECT 13.280 51.175 13.630 53.335 ;
        RECT 14.110 51.175 14.460 53.335 ;
        RECT 14.940 51.175 15.290 53.335 ;
        RECT 15.770 51.175 16.120 53.335 ;
        RECT 16.600 51.175 16.950 53.335 ;
        RECT 17.430 51.175 17.780 53.335 ;
        RECT 18.260 51.175 18.610 53.335 ;
        RECT 19.090 51.175 19.440 53.335 ;
        RECT 0.000 17.175 0.350 19.335 ;
        RECT 0.830 17.175 1.180 19.335 ;
        RECT 1.660 17.175 2.010 19.335 ;
        RECT 2.490 17.175 2.840 19.335 ;
        RECT 3.320 17.175 3.670 19.335 ;
        RECT 4.150 17.175 4.500 19.335 ;
        RECT 4.980 17.175 5.330 19.335 ;
        RECT 5.810 17.175 6.160 19.335 ;
        RECT 6.640 17.175 6.990 19.335 ;
        RECT 7.470 17.175 7.820 19.335 ;
        RECT 8.300 17.175 8.650 19.335 ;
        RECT 9.130 17.175 9.480 19.335 ;
        RECT 9.960 17.175 10.310 19.335 ;
        RECT 10.790 17.175 11.140 19.335 ;
        RECT 11.620 17.175 11.970 19.335 ;
        RECT 12.450 17.175 12.800 19.335 ;
        RECT 13.280 17.175 13.630 19.335 ;
        RECT 14.110 17.175 14.460 19.335 ;
        RECT 14.940 17.175 15.290 19.335 ;
        RECT 15.770 17.175 16.120 19.335 ;
        RECT 16.600 17.175 16.950 19.335 ;
        RECT 17.430 17.175 17.780 19.335 ;
        RECT 18.260 17.175 18.610 19.335 ;
        RECT 19.090 17.175 19.440 19.335 ;
        RECT 0.000 14.740 0.350 16.900 ;
        RECT 0.830 14.740 1.180 16.900 ;
        RECT 1.660 14.740 2.010 16.900 ;
        RECT 2.490 14.740 2.840 16.900 ;
        RECT 3.610 16.135 4.610 16.305 ;
        RECT 4.970 16.240 5.180 16.610 ;
        RECT 5.490 16.135 6.490 16.305 ;
        RECT 6.850 16.240 7.060 16.610 ;
        RECT 7.370 16.135 8.370 16.305 ;
        RECT 8.730 16.240 8.940 16.610 ;
        RECT 9.250 16.135 10.250 16.305 ;
        RECT 10.610 16.240 10.820 16.610 ;
        RECT 11.130 16.135 12.130 16.305 ;
        RECT 12.490 16.240 12.700 16.610 ;
        RECT 13.010 16.135 14.010 16.305 ;
        RECT 3.380 11.880 3.550 15.920 ;
        RECT 4.670 11.880 4.840 15.920 ;
        RECT 5.260 11.880 5.430 15.920 ;
        RECT 6.550 11.880 6.720 15.920 ;
        RECT 7.140 11.880 7.310 15.920 ;
        RECT 8.430 11.880 8.600 15.920 ;
        RECT 9.020 11.880 9.190 15.920 ;
        RECT 10.310 11.880 10.480 15.920 ;
        RECT 10.900 11.880 11.070 15.920 ;
        RECT 12.190 11.880 12.360 15.920 ;
        RECT 12.780 11.880 12.950 15.920 ;
        RECT 14.070 11.880 14.240 15.920 ;
        RECT 3.610 11.495 4.610 11.665 ;
        RECT 5.490 11.495 6.490 11.665 ;
        RECT 7.370 11.495 8.370 11.665 ;
        RECT 9.250 11.495 10.250 11.665 ;
        RECT 11.130 11.495 12.130 11.665 ;
        RECT 13.010 11.495 14.010 11.665 ;
        RECT 3.610 10.955 4.610 11.125 ;
        RECT 5.490 10.955 6.490 11.125 ;
        RECT 7.370 10.955 8.370 11.125 ;
        RECT 9.250 10.955 10.250 11.125 ;
        RECT 11.130 10.955 12.130 11.125 ;
        RECT 13.010 10.955 14.010 11.125 ;
        RECT 0.000 6.490 0.350 8.650 ;
        RECT 0.830 6.490 1.180 8.650 ;
        RECT 1.660 6.490 2.010 8.650 ;
        RECT 2.490 6.490 2.840 8.650 ;
        RECT 3.380 6.700 3.550 10.740 ;
        RECT 4.670 6.700 4.840 10.740 ;
        RECT 5.260 6.700 5.430 10.740 ;
        RECT 6.550 6.700 6.720 10.740 ;
        RECT 7.140 6.700 7.310 10.740 ;
        RECT 8.430 6.700 8.600 10.740 ;
        RECT 9.020 6.700 9.190 10.740 ;
        RECT 10.310 6.700 10.480 10.740 ;
        RECT 10.900 6.700 11.070 10.740 ;
        RECT 12.190 6.700 12.360 10.740 ;
        RECT 12.780 6.700 12.950 10.740 ;
        RECT 14.070 6.700 14.240 10.740 ;
        RECT 3.610 6.315 4.610 6.485 ;
        RECT 5.490 6.315 6.490 6.485 ;
        RECT 7.370 6.315 8.370 6.485 ;
        RECT 9.250 6.315 10.250 6.485 ;
        RECT 11.130 6.315 12.130 6.485 ;
        RECT 13.010 6.315 14.010 6.485 ;
        RECT 1.730 5.760 2.730 5.930 ;
        RECT 3.610 5.760 4.610 5.930 ;
        RECT 5.490 5.760 6.490 5.930 ;
        RECT 7.370 5.760 8.370 5.930 ;
        RECT 9.250 5.760 10.250 5.930 ;
        RECT 11.130 5.760 12.130 5.930 ;
        RECT 13.010 5.760 14.010 5.930 ;
        RECT 0.030 4.810 0.240 5.180 ;
        RECT 0.030 3.525 0.240 3.895 ;
        RECT 1.500 3.550 1.670 5.590 ;
        RECT 2.790 3.550 2.960 5.590 ;
        RECT 3.380 3.550 3.550 5.590 ;
        RECT 4.670 3.550 4.840 5.590 ;
        RECT 5.260 3.550 5.430 5.590 ;
        RECT 6.550 3.550 6.720 5.590 ;
        RECT 7.140 3.550 7.310 5.590 ;
        RECT 8.430 3.550 8.600 5.590 ;
        RECT 9.020 3.550 9.190 5.590 ;
        RECT 10.310 3.550 10.480 5.590 ;
        RECT 10.900 3.550 11.070 5.590 ;
        RECT 12.190 3.550 12.360 5.590 ;
        RECT 12.780 3.550 12.950 5.590 ;
        RECT 14.070 3.550 14.240 5.590 ;
        RECT 1.730 3.210 2.730 3.380 ;
        RECT 3.610 3.210 4.610 3.380 ;
        RECT 5.490 3.210 6.490 3.380 ;
        RECT 7.370 3.210 8.370 3.380 ;
        RECT 9.250 3.210 10.250 3.380 ;
        RECT 11.130 3.210 12.130 3.380 ;
        RECT 13.010 3.210 14.010 3.380 ;
        RECT 1.730 2.670 2.730 2.840 ;
        RECT 3.610 2.670 4.610 2.840 ;
        RECT 5.490 2.670 6.490 2.840 ;
        RECT 7.370 2.670 8.370 2.840 ;
        RECT 9.250 2.670 10.250 2.840 ;
        RECT 11.130 2.670 12.130 2.840 ;
        RECT 13.010 2.670 14.010 2.840 ;
        RECT 0.030 2.240 0.240 2.610 ;
        RECT 0.030 0.950 0.240 1.320 ;
        RECT 1.500 0.460 1.670 2.500 ;
        RECT 2.790 0.460 2.960 2.500 ;
        RECT 3.380 0.460 3.550 2.500 ;
        RECT 4.670 0.460 4.840 2.500 ;
        RECT 5.260 0.460 5.430 2.500 ;
        RECT 6.550 0.460 6.720 2.500 ;
        RECT 7.140 0.460 7.310 2.500 ;
        RECT 8.430 0.460 8.600 2.500 ;
        RECT 9.020 0.460 9.190 2.500 ;
        RECT 10.310 0.460 10.480 2.500 ;
        RECT 10.900 0.460 11.070 2.500 ;
        RECT 12.190 0.460 12.360 2.500 ;
        RECT 12.780 0.460 12.950 2.500 ;
        RECT 14.070 0.460 14.240 2.500 ;
        RECT 1.730 0.120 2.730 0.290 ;
        RECT 3.610 0.120 4.610 0.290 ;
        RECT 5.490 0.120 6.490 0.290 ;
        RECT 7.370 0.120 8.370 0.290 ;
        RECT 9.250 0.120 10.250 0.290 ;
        RECT 11.130 0.120 12.130 0.290 ;
        RECT 13.010 0.120 14.010 0.290 ;
        RECT 20.325 -1.320 20.495 53.960 ;
        RECT -2.305 -1.490 20.495 -1.320 ;
      LAYER met1 ;
        RECT 0.000 51.175 1.180 53.335 ;
        RECT 1.660 51.175 2.840 53.335 ;
        RECT 3.320 51.175 4.500 53.335 ;
        RECT 4.980 51.175 6.160 53.335 ;
        RECT 6.640 51.175 7.820 53.335 ;
        RECT 8.300 51.175 9.480 53.335 ;
        RECT 9.960 51.175 11.140 53.335 ;
        RECT 11.620 51.175 12.800 53.335 ;
        RECT 13.280 51.175 14.460 53.335 ;
        RECT 14.940 51.175 16.120 53.335 ;
        RECT 16.600 51.175 17.780 53.335 ;
        RECT 18.260 51.175 19.440 53.335 ;
        RECT 0.000 17.175 0.350 19.335 ;
        RECT 0.830 17.175 2.010 19.335 ;
        RECT 2.490 17.175 3.670 19.335 ;
        RECT 4.150 17.175 5.330 19.335 ;
        RECT 5.810 17.175 6.990 19.335 ;
        RECT 7.470 17.175 8.650 19.335 ;
        RECT 9.130 17.175 10.310 19.335 ;
        RECT 10.790 17.175 11.970 19.335 ;
        RECT 12.450 17.175 13.630 19.335 ;
        RECT 14.110 17.175 15.290 19.335 ;
        RECT 15.770 17.175 16.950 19.335 ;
        RECT 17.430 17.175 18.610 19.335 ;
        RECT 19.090 17.175 19.440 19.335 ;
        RECT 0.000 14.740 1.190 16.900 ;
        RECT 1.660 14.740 2.850 16.900 ;
        RECT 4.910 16.645 12.760 16.835 ;
        RECT 3.630 16.330 4.590 16.335 ;
        RECT 3.350 16.105 4.590 16.330 ;
        RECT 4.910 16.260 5.240 16.645 ;
        RECT 5.510 16.105 6.470 16.335 ;
        RECT 6.790 16.260 7.120 16.645 ;
        RECT 7.390 16.330 8.350 16.430 ;
        RECT 7.260 16.120 8.350 16.330 ;
        RECT 8.670 16.260 9.000 16.645 ;
        RECT 3.350 15.670 4.210 16.105 ;
        RECT 3.350 12.145 3.580 15.670 ;
        RECT 3.265 12.140 3.580 12.145 ;
        RECT 4.015 12.140 4.205 15.670 ;
        RECT 4.350 15.310 4.950 15.910 ;
        RECT 3.265 11.700 4.205 12.140 ;
        RECT 4.640 12.155 4.870 15.310 ;
        RECT 4.640 11.900 4.965 12.155 ;
        RECT 5.230 12.140 5.460 15.900 ;
        RECT 3.265 10.920 4.610 11.700 ;
        RECT 3.265 10.480 4.205 10.920 ;
        RECT 4.775 10.720 4.965 11.900 ;
        RECT 3.265 10.475 3.580 10.480 ;
        RECT 0.000 6.460 0.350 8.680 ;
        RECT 0.830 6.490 2.020 8.650 ;
        RECT 2.540 5.960 2.790 8.625 ;
        RECT 3.350 7.260 3.580 10.475 ;
        RECT 3.160 6.950 3.770 7.260 ;
        RECT 4.015 6.950 4.205 10.480 ;
        RECT 4.640 10.495 4.965 10.720 ;
        RECT 5.145 11.900 5.460 12.140 ;
        RECT 5.145 10.720 5.335 11.900 ;
        RECT 5.895 11.700 6.085 16.105 ;
        RECT 7.140 16.100 8.350 16.120 ;
        RECT 9.270 16.100 10.230 16.430 ;
        RECT 10.550 16.260 10.880 16.645 ;
        RECT 6.240 15.310 6.840 15.910 ;
        RECT 7.140 15.900 7.965 16.100 ;
        RECT 7.110 15.670 7.965 15.900 ;
        RECT 6.520 12.140 6.750 15.310 ;
        RECT 7.110 12.150 7.340 15.670 ;
        RECT 7.775 12.150 7.965 15.670 ;
        RECT 7.030 12.145 7.965 12.150 ;
        RECT 6.520 11.900 6.845 12.140 ;
        RECT 5.490 10.920 6.490 11.700 ;
        RECT 5.145 10.515 5.460 10.720 ;
        RECT 3.160 6.660 4.210 6.950 ;
        RECT 4.640 6.720 4.870 10.495 ;
        RECT 5.230 7.260 5.460 10.515 ;
        RECT 5.040 6.660 5.650 7.260 ;
        RECT 3.380 6.515 4.210 6.660 ;
        RECT 5.895 6.515 6.085 10.920 ;
        RECT 6.655 10.720 6.845 11.900 ;
        RECT 6.520 10.485 6.845 10.720 ;
        RECT 7.025 11.700 7.965 12.145 ;
        RECT 8.400 15.360 9.220 15.900 ;
        RECT 8.400 12.140 8.630 15.360 ;
        RECT 8.990 12.140 9.220 15.360 ;
        RECT 8.400 11.900 9.220 12.140 ;
        RECT 7.025 10.920 8.350 11.700 ;
        RECT 7.025 10.490 7.970 10.920 ;
        RECT 8.525 10.720 9.085 11.900 ;
        RECT 9.655 11.700 9.845 16.100 ;
        RECT 11.150 16.060 12.110 16.380 ;
        RECT 12.430 16.260 12.760 16.645 ;
        RECT 13.030 16.060 13.990 16.380 ;
        RECT 10.280 12.140 10.510 15.900 ;
        RECT 10.870 12.145 11.100 15.900 ;
        RECT 10.280 11.900 10.615 12.140 ;
        RECT 9.270 10.920 10.230 11.700 ;
        RECT 7.025 10.485 7.965 10.490 ;
        RECT 6.520 6.720 6.750 10.485 ;
        RECT 7.030 10.480 7.965 10.485 ;
        RECT 7.110 6.960 7.340 10.480 ;
        RECT 7.015 6.950 7.340 6.960 ;
        RECT 7.775 6.950 7.965 10.480 ;
        RECT 8.400 10.470 9.220 10.720 ;
        RECT 8.400 6.960 8.630 10.470 ;
        RECT 8.990 6.960 9.220 10.470 ;
        RECT 7.015 6.515 7.970 6.950 ;
        RECT 8.400 6.770 9.220 6.960 ;
        RECT 8.400 6.720 8.630 6.770 ;
        RECT 8.990 6.720 9.220 6.770 ;
        RECT 9.655 6.515 9.845 10.920 ;
        RECT 10.425 10.720 10.615 11.900 ;
        RECT 10.280 10.485 10.615 10.720 ;
        RECT 10.785 11.900 11.100 12.145 ;
        RECT 10.785 10.720 10.975 11.900 ;
        RECT 11.535 11.695 11.725 16.060 ;
        RECT 12.160 15.850 12.390 15.900 ;
        RECT 12.750 15.850 12.980 15.900 ;
        RECT 12.160 15.660 12.980 15.850 ;
        RECT 12.160 12.135 12.390 15.660 ;
        RECT 12.750 12.140 12.980 15.660 ;
        RECT 12.635 12.135 12.980 12.140 ;
        RECT 12.160 11.900 12.980 12.135 ;
        RECT 11.150 11.465 12.110 11.695 ;
        RECT 11.160 11.155 12.100 11.465 ;
        RECT 12.285 11.400 12.825 11.900 ;
        RECT 13.415 11.695 13.605 16.060 ;
        RECT 14.040 12.140 14.270 15.900 ;
        RECT 14.040 11.900 14.355 12.140 ;
        RECT 13.030 11.465 13.990 11.695 ;
        RECT 12.285 11.210 12.835 11.400 ;
        RECT 11.150 10.925 12.110 11.155 ;
        RECT 10.785 10.485 11.100 10.720 ;
        RECT 10.280 7.330 10.510 10.485 ;
        RECT 10.000 6.730 10.610 7.330 ;
        RECT 10.870 6.965 11.100 10.485 ;
        RECT 10.280 6.720 10.610 6.730 ;
        RECT 3.380 6.320 4.590 6.515 ;
        RECT 3.630 6.285 4.590 6.320 ;
        RECT 5.510 6.285 6.470 6.515 ;
        RECT 7.015 6.510 8.350 6.515 ;
        RECT 9.270 6.510 10.230 6.515 ;
        RECT 7.015 6.280 10.230 6.510 ;
        RECT 1.470 5.730 6.490 5.960 ;
        RECT 1.470 5.340 2.330 5.730 ;
        RECT 0.000 5.090 0.270 5.180 ;
        RECT 0.000 4.900 1.225 5.090 ;
        RECT 0.000 4.800 0.270 4.900 ;
        RECT 0.040 4.765 0.230 4.800 ;
        RECT 0.000 3.805 0.270 3.895 ;
        RECT 1.035 3.805 1.225 4.900 ;
        RECT 1.470 3.820 1.700 5.340 ;
        RECT 2.135 3.820 2.330 5.340 ;
        RECT 1.380 3.815 2.330 3.820 ;
        RECT 0.000 3.615 1.225 3.805 ;
        RECT 0.000 3.515 0.270 3.615 ;
        RECT 0.040 3.485 0.230 3.515 ;
        RECT 0.000 2.520 0.270 2.610 ;
        RECT 1.035 2.520 1.225 3.615 ;
        RECT 0.000 2.330 1.225 2.520 ;
        RECT 0.000 2.230 0.270 2.330 ;
        RECT 0.040 2.200 0.230 2.230 ;
        RECT 0.000 1.230 0.270 1.320 ;
        RECT 1.035 1.230 1.225 2.330 ;
        RECT 1.375 3.410 2.330 3.815 ;
        RECT 2.760 3.815 2.990 5.570 ;
        RECT 3.350 5.560 3.580 5.570 ;
        RECT 3.160 4.960 3.760 5.560 ;
        RECT 2.760 3.570 3.085 3.815 ;
        RECT 3.350 3.810 3.580 4.960 ;
        RECT 1.375 2.640 2.730 3.410 ;
        RECT 1.375 2.250 2.330 2.640 ;
        RECT 2.895 2.480 3.085 3.570 ;
        RECT 1.375 2.240 1.700 2.250 ;
        RECT 0.000 1.040 1.225 1.230 ;
        RECT 0.000 0.940 0.270 1.040 ;
        RECT 1.000 0.990 1.225 1.040 ;
        RECT 0.040 0.910 0.230 0.940 ;
        RECT 1.000 0.670 1.260 0.990 ;
        RECT 1.470 0.720 1.700 2.240 ;
        RECT 2.135 0.720 2.330 2.250 ;
        RECT 2.760 2.225 3.085 2.480 ;
        RECT 3.265 3.570 3.580 3.810 ;
        RECT 3.265 2.480 3.455 3.570 ;
        RECT 4.015 3.410 4.205 5.730 ;
        RECT 4.640 3.810 4.870 5.570 ;
        RECT 5.230 5.560 5.460 5.570 ;
        RECT 5.040 4.960 5.640 5.560 ;
        RECT 5.230 3.815 5.460 4.960 ;
        RECT 4.640 3.570 4.965 3.810 ;
        RECT 3.610 2.640 4.610 3.410 ;
        RECT 3.265 2.225 3.580 2.480 ;
        RECT 2.760 1.080 2.990 2.225 ;
        RECT 1.470 0.320 2.330 0.720 ;
        RECT 2.470 0.480 3.070 1.080 ;
        RECT 3.350 0.480 3.580 2.225 ;
        RECT 4.015 0.320 4.205 2.640 ;
        RECT 4.775 2.480 4.965 3.570 ;
        RECT 4.640 2.225 4.965 2.480 ;
        RECT 5.145 3.570 5.460 3.815 ;
        RECT 5.145 2.480 5.335 3.570 ;
        RECT 5.895 3.410 6.085 5.730 ;
        RECT 7.015 5.570 7.205 6.280 ;
        RECT 7.390 5.730 8.350 5.960 ;
        RECT 9.270 5.730 10.230 5.960 ;
        RECT 6.520 3.810 6.750 5.570 ;
        RECT 7.015 5.325 7.340 5.570 ;
        RECT 7.110 3.815 7.340 5.325 ;
        RECT 6.520 3.570 6.835 3.810 ;
        RECT 5.490 2.640 6.490 3.410 ;
        RECT 5.145 2.235 5.460 2.480 ;
        RECT 4.640 1.080 4.870 2.225 ;
        RECT 4.350 0.480 4.950 1.080 ;
        RECT 5.230 0.480 5.460 2.235 ;
        RECT 5.895 0.320 6.085 2.640 ;
        RECT 6.645 2.480 6.835 3.570 ;
        RECT 6.520 2.235 6.835 2.480 ;
        RECT 7.025 3.570 7.340 3.815 ;
        RECT 7.025 2.480 7.215 3.570 ;
        RECT 7.775 3.410 7.965 5.730 ;
        RECT 8.400 5.520 8.630 5.570 ;
        RECT 8.990 5.520 9.220 5.570 ;
        RECT 8.400 5.330 9.220 5.520 ;
        RECT 8.400 3.810 8.630 5.330 ;
        RECT 8.990 3.810 9.220 5.330 ;
        RECT 8.400 3.570 9.220 3.810 ;
        RECT 7.390 2.640 8.350 3.410 ;
        RECT 7.025 2.240 7.340 2.480 ;
        RECT 6.520 1.080 6.750 2.235 ;
        RECT 6.230 0.480 6.830 1.080 ;
        RECT 7.110 0.480 7.340 2.240 ;
        RECT 7.775 0.320 7.965 2.640 ;
        RECT 8.525 2.480 9.085 3.570 ;
        RECT 9.655 3.410 9.845 5.730 ;
        RECT 10.420 5.570 10.610 6.720 ;
        RECT 10.280 5.560 10.610 5.570 ;
        RECT 10.000 4.960 10.610 5.560 ;
        RECT 10.785 6.720 11.100 6.965 ;
        RECT 10.785 5.960 10.975 6.720 ;
        RECT 11.535 6.515 11.725 10.925 ;
        RECT 12.285 10.720 12.825 11.210 ;
        RECT 13.090 11.155 13.930 11.465 ;
        RECT 13.030 10.925 13.990 11.155 ;
        RECT 12.160 10.480 12.980 10.720 ;
        RECT 12.160 6.960 12.390 10.480 ;
        RECT 12.635 10.475 12.980 10.480 ;
        RECT 12.750 6.960 12.980 10.475 ;
        RECT 12.160 6.770 12.980 6.960 ;
        RECT 12.160 6.720 12.390 6.770 ;
        RECT 12.750 6.720 12.980 6.770 ;
        RECT 13.415 6.515 13.605 10.925 ;
        RECT 14.165 10.720 14.355 11.900 ;
        RECT 14.040 10.475 14.355 10.720 ;
        RECT 14.040 7.320 14.270 10.475 ;
        RECT 13.810 6.720 14.410 7.320 ;
        RECT 11.150 6.285 12.110 6.515 ;
        RECT 13.030 6.285 13.990 6.515 ;
        RECT 10.785 5.940 12.110 5.960 ;
        RECT 13.030 5.940 13.990 5.960 ;
        RECT 10.785 5.750 13.990 5.940 ;
        RECT 10.785 5.730 12.110 5.750 ;
        RECT 13.030 5.730 13.990 5.750 ;
        RECT 10.785 5.325 11.730 5.730 ;
        RECT 10.790 5.320 11.730 5.325 ;
        RECT 12.160 5.520 12.390 5.570 ;
        RECT 12.750 5.520 12.980 5.570 ;
        RECT 12.160 5.330 12.980 5.520 ;
        RECT 10.280 3.810 10.510 4.960 ;
        RECT 10.870 3.810 11.100 5.320 ;
        RECT 11.535 3.810 11.725 5.320 ;
        RECT 10.280 3.570 10.595 3.810 ;
        RECT 9.270 2.640 10.230 3.410 ;
        RECT 8.400 2.240 9.220 2.480 ;
        RECT 8.400 0.720 8.630 2.240 ;
        RECT 8.990 0.720 9.220 2.240 ;
        RECT 8.400 0.530 9.220 0.720 ;
        RECT 8.400 0.480 8.630 0.530 ;
        RECT 8.990 0.480 9.220 0.530 ;
        RECT 9.655 0.320 9.845 2.640 ;
        RECT 10.405 2.480 10.595 3.570 ;
        RECT 10.280 2.225 10.595 2.480 ;
        RECT 10.775 3.420 11.725 3.810 ;
        RECT 12.160 3.810 12.390 5.330 ;
        RECT 12.750 3.810 12.980 5.330 ;
        RECT 12.160 3.570 12.980 3.810 ;
        RECT 10.775 2.640 12.110 3.420 ;
        RECT 10.775 2.240 11.725 2.640 ;
        RECT 12.295 2.480 12.860 3.570 ;
        RECT 13.415 3.410 13.605 5.730 ;
        RECT 14.215 5.570 14.410 6.720 ;
        RECT 13.810 4.960 14.410 5.570 ;
        RECT 14.040 3.810 14.270 4.960 ;
        RECT 14.040 3.570 14.355 3.810 ;
        RECT 13.030 2.640 13.990 3.410 ;
        RECT 10.775 2.235 11.100 2.240 ;
        RECT 10.280 0.480 10.510 2.225 ;
        RECT 10.870 0.710 11.100 2.235 ;
        RECT 11.535 0.710 11.725 2.240 ;
        RECT 12.160 2.230 12.980 2.480 ;
        RECT 12.160 1.110 12.390 2.230 ;
        RECT 12.750 1.110 12.980 2.230 ;
        RECT 10.870 0.480 11.730 0.710 ;
        RECT 12.160 0.510 12.980 1.110 ;
        RECT 12.160 0.480 12.390 0.510 ;
        RECT 12.750 0.480 12.980 0.510 ;
        RECT 10.890 0.360 11.730 0.480 ;
        RECT 13.415 0.360 13.605 2.640 ;
        RECT 14.165 2.480 14.355 3.570 ;
        RECT 14.040 2.245 14.355 2.480 ;
        RECT 14.040 0.480 14.270 2.245 ;
        RECT 10.890 0.320 12.080 0.360 ;
        RECT 13.060 0.320 13.960 0.360 ;
        RECT 1.470 0.090 2.730 0.320 ;
        RECT 1.730 0.000 2.730 0.090 ;
        RECT 3.610 0.000 4.610 0.320 ;
        RECT 5.490 0.000 6.490 0.320 ;
        RECT 7.390 0.090 8.350 0.320 ;
        RECT 9.270 0.090 10.230 0.320 ;
        RECT 10.890 0.115 12.110 0.320 ;
        RECT 11.150 0.090 12.110 0.115 ;
        RECT 13.030 0.090 13.990 0.320 ;
        RECT 11.180 0.040 12.080 0.090 ;
        RECT 13.060 0.040 13.960 0.090 ;
      LAYER met2 ;
        RECT 0.000 17.175 0.350 19.335 ;
        RECT 5.900 17.755 6.900 18.755 ;
        RECT 12.510 17.785 13.570 18.725 ;
        RECT 0.055 16.980 0.295 17.175 ;
        RECT 12.915 16.980 13.160 17.785 ;
        RECT 19.090 17.175 19.440 19.335 ;
        RECT 19.140 16.980 19.380 17.175 ;
        RECT 0.055 16.740 11.750 16.980 ;
        RECT 4.915 16.300 5.235 16.560 ;
        RECT 4.950 15.910 5.200 16.300 ;
        RECT 7.390 16.110 10.230 16.430 ;
        RECT 11.510 16.380 11.750 16.740 ;
        RECT 12.915 16.735 13.635 16.980 ;
        RECT 14.400 16.740 19.380 16.980 ;
        RECT 13.390 16.380 13.630 16.735 ;
        RECT 11.150 16.060 12.110 16.380 ;
        RECT 13.030 16.060 13.990 16.380 ;
        RECT 4.350 15.750 5.350 15.910 ;
        RECT 6.240 15.750 7.240 15.910 ;
        RECT 8.300 15.750 9.300 15.900 ;
        RECT 0.050 15.510 9.300 15.750 ;
        RECT 0.050 8.680 0.290 15.510 ;
        RECT 4.350 14.910 5.350 15.510 ;
        RECT 6.240 14.910 7.240 15.510 ;
        RECT 8.300 14.900 9.300 15.510 ;
        RECT 6.770 12.410 12.675 12.650 ;
        RECT 3.610 11.435 4.610 11.700 ;
        RECT 5.490 11.435 6.490 11.700 ;
        RECT 3.610 11.185 6.490 11.435 ;
        RECT 3.610 10.920 4.610 11.185 ;
        RECT 5.490 10.920 6.490 11.185 ;
        RECT 0.000 6.460 0.350 8.680 ;
        RECT 3.160 6.660 3.770 7.260 ;
        RECT 5.040 7.080 5.650 7.260 ;
        RECT 6.770 7.080 7.010 12.410 ;
        RECT 12.435 12.130 12.675 12.410 ;
        RECT 7.390 11.435 8.350 11.700 ;
        RECT 9.270 11.435 10.230 11.700 ;
        RECT 7.390 11.185 10.230 11.435 ;
        RECT 7.390 10.920 8.350 11.185 ;
        RECT 9.270 10.920 10.230 11.185 ;
        RECT 11.160 10.930 12.100 11.690 ;
        RECT 11.510 9.270 11.750 10.930 ;
        RECT 12.290 10.490 12.820 12.130 ;
        RECT 13.030 10.930 13.990 11.690 ;
        RECT 5.040 6.840 7.010 7.080 ;
        RECT 7.740 9.030 11.750 9.270 ;
        RECT 5.040 6.660 5.650 6.840 ;
        RECT 0.050 6.140 0.300 6.460 ;
        RECT 0.000 5.140 1.000 6.140 ;
        RECT 3.335 5.560 3.585 6.660 ;
        RECT 7.740 6.230 7.980 9.030 ;
        RECT 13.390 8.220 13.630 10.930 ;
        RECT 4.560 5.990 7.980 6.230 ;
        RECT 3.160 4.960 3.760 5.560 ;
        RECT 0.000 4.580 1.000 4.850 ;
        RECT 4.560 4.580 4.800 5.990 ;
        RECT 5.040 5.390 5.640 5.560 ;
        RECT 5.040 5.150 7.050 5.390 ;
        RECT 5.040 4.960 5.640 5.150 ;
        RECT 0.000 4.340 4.800 4.580 ;
        RECT 0.000 3.850 1.000 4.340 ;
        RECT 0.000 3.030 1.000 3.570 ;
        RECT 1.730 3.150 2.730 3.410 ;
        RECT 3.610 3.150 4.610 3.410 ;
        RECT 5.490 3.150 6.490 3.410 ;
        RECT 0.000 2.790 1.440 3.030 ;
        RECT 0.000 2.570 1.000 2.790 ;
        RECT 0.000 1.635 1.000 2.270 ;
        RECT 1.200 2.070 1.440 2.790 ;
        RECT 1.730 2.900 6.490 3.150 ;
        RECT 1.730 2.640 2.730 2.900 ;
        RECT 3.610 2.640 4.610 2.900 ;
        RECT 5.490 2.640 6.490 2.900 ;
        RECT 6.810 2.490 7.050 5.150 ;
        RECT 7.740 3.410 7.980 5.990 ;
        RECT 9.620 7.980 13.630 8.220 ;
        RECT 7.390 2.640 8.350 3.410 ;
        RECT 8.525 2.490 9.085 3.810 ;
        RECT 9.620 3.410 9.860 7.980 ;
        RECT 14.400 7.730 14.640 16.740 ;
        RECT 10.000 6.730 10.610 7.330 ;
        RECT 13.640 6.730 14.640 7.730 ;
        RECT 10.180 6.245 10.430 6.730 ;
        RECT 13.990 6.245 14.240 6.730 ;
        RECT 10.180 5.995 14.240 6.245 ;
        RECT 10.180 5.560 10.430 5.995 ;
        RECT 13.990 5.570 14.240 5.995 ;
        RECT 10.000 4.960 10.610 5.560 ;
        RECT 13.810 4.960 14.410 5.570 ;
        RECT 10.180 4.055 10.430 4.960 ;
        RECT 10.180 3.805 10.665 4.055 ;
        RECT 9.270 2.640 10.230 3.410 ;
        RECT 6.810 2.250 9.085 2.490 ;
        RECT 9.630 2.070 9.870 2.640 ;
        RECT 1.200 1.830 9.870 2.070 ;
        RECT 10.415 1.635 10.665 3.805 ;
        RECT 11.140 3.150 12.110 3.420 ;
        RECT 13.030 3.150 13.990 3.410 ;
        RECT 11.140 2.900 13.990 3.150 ;
        RECT 11.140 2.640 12.110 2.900 ;
        RECT 13.030 2.640 13.990 2.900 ;
        RECT 0.000 1.385 10.665 1.635 ;
        RECT 0.000 1.270 1.000 1.385 ;
        RECT 0.000 0.960 1.000 1.000 ;
        RECT 0.000 0.930 1.290 0.960 ;
        RECT 2.100 0.930 3.420 1.230 ;
        RECT 3.980 0.930 5.300 1.240 ;
        RECT 5.860 0.930 7.180 1.240 ;
        RECT 11.900 0.930 13.220 1.260 ;
        RECT 0.000 0.690 13.220 0.930 ;
        RECT 0.000 0.000 1.000 0.690 ;
        RECT 2.100 0.470 3.420 0.690 ;
        RECT 3.980 0.480 5.300 0.690 ;
        RECT 5.860 0.480 7.180 0.690 ;
        RECT 11.900 0.500 13.220 0.690 ;
        RECT 11.150 0.330 12.130 0.360 ;
        RECT 13.010 0.330 14.000 0.360 ;
        RECT 1.730 0.285 2.730 0.320 ;
        RECT 3.610 0.285 4.610 0.320 ;
        RECT 5.490 0.285 6.490 0.320 ;
        RECT 1.730 0.035 6.490 0.285 ;
        RECT 11.150 0.080 14.000 0.330 ;
        RECT 11.150 0.040 12.130 0.080 ;
        RECT 13.010 0.040 14.000 0.080 ;
        RECT 1.730 0.000 2.730 0.035 ;
        RECT 3.610 0.000 4.610 0.035 ;
        RECT 5.490 0.000 6.490 0.035 ;
      LAYER met3 ;
        RECT 4.350 11.820 5.350 15.910 ;
        RECT 6.240 11.820 7.240 15.910 ;
        RECT 8.300 11.820 9.300 15.900 ;
        RECT 3.260 10.820 14.350 11.820 ;
        RECT 0.000 5.140 1.000 6.140 ;
        RECT 1.380 2.570 14.350 3.570 ;
        RECT 2.260 1.230 3.260 2.570 ;
        RECT 4.140 1.240 5.140 2.570 ;
        RECT 6.020 1.240 7.020 2.570 ;
        RECT 12.060 1.260 13.060 2.570 ;
        RECT 0.000 0.000 1.000 1.000 ;
        RECT 2.100 0.470 3.420 1.230 ;
        RECT 3.980 0.480 5.300 1.240 ;
        RECT 5.860 0.480 7.180 1.240 ;
        RECT 11.900 0.500 13.220 1.260 ;
        RECT 2.260 0.350 3.260 0.470 ;
        RECT 4.140 0.360 5.140 0.480 ;
        RECT 6.020 0.360 7.020 0.480 ;
        RECT 12.060 0.380 13.060 0.500 ;
  END
END hybrid_dnwell
END LIBRARY

