magic
tech sky130A
magscale 1 2
timestamp 1727607728
<< dnwell >>
rect -606 4500 3302 6733
rect -606 -335 3302 3240
<< nwell >>
rect -686 6527 3382 6813
rect -686 4706 -400 6527
rect 3096 4706 3382 6527
rect -686 4420 3382 4706
rect -686 3034 3382 3320
rect -686 -129 -400 3034
rect 3096 -129 3382 3034
rect -686 -415 3382 -129
<< nsubdiff >>
rect -649 6756 3345 6776
rect -649 6722 -569 6756
rect 3265 6722 3345 6756
rect -649 6702 3345 6722
rect -649 6696 -575 6702
rect -649 4537 -629 6696
rect -595 4537 -575 6696
rect -649 4531 -575 4537
rect 3271 6696 3345 6702
rect 3271 4537 3291 6696
rect 3325 4537 3345 6696
rect 3271 4531 3345 4537
rect -649 4511 3345 4531
rect -649 4477 -569 4511
rect 3265 4477 3345 4511
rect -649 4457 3345 4477
rect -649 3263 3345 3283
rect -649 3229 -569 3263
rect 3265 3229 3345 3263
rect -649 3209 3345 3229
rect -649 3203 -575 3209
rect -649 -298 -629 3203
rect -595 -298 -575 3203
rect -649 -304 -575 -298
rect 3271 3203 3345 3209
rect 3271 -298 3291 3203
rect 3325 -298 3345 3203
rect 3271 -304 3345 -298
rect -649 -324 3345 -304
rect -649 -358 -569 -324
rect 3265 -358 3345 -324
rect -649 -378 3345 -358
<< nsubdiffcont >>
rect -569 6722 3265 6756
rect -629 4537 -595 6696
rect 3291 4537 3325 6696
rect -569 4477 3265 4511
rect -569 3229 3265 3263
rect -629 -298 -595 3203
rect 3291 -298 3325 3203
rect -569 -358 3265 -324
<< locali >>
rect -629 6722 -569 6756
rect 3265 6722 3325 6756
rect -629 6696 -595 6722
rect -629 4511 -595 4537
rect 3291 6696 3325 6722
rect 3291 4511 3325 4537
rect -629 4477 -569 4511
rect 3265 4477 3325 4511
rect -629 3229 -569 3263
rect 3265 3229 3325 3263
rect -629 3203 -595 3229
rect -629 -324 -595 -298
rect 3291 3203 3325 3229
rect 3291 -324 3325 -298
rect -629 -358 -569 -324
rect 3265 -358 3325 -324
use shifters_split  shifters_split_0
timestamp 1727607728
transform 1 0 60 0 1 0
box -60 0 2636 6127
<< end >>
