magic
tech sky130A
magscale 1 2
timestamp 1727641294
<< nwell >>
rect -48 954 524 2076
<< pwell >>
rect -48 0 527 905
<< mvnmos >>
rect 188 561 288 691
rect 188 213 288 343
<< mvpmos >>
rect 188 1633 288 1833
rect 188 1197 288 1397
<< mvndiff >>
rect 130 679 188 691
rect 130 573 142 679
rect 176 573 188 679
rect 130 561 188 573
rect 288 679 346 691
rect 288 573 300 679
rect 334 573 346 679
rect 288 561 346 573
rect 130 331 188 343
rect 130 225 142 331
rect 176 225 188 331
rect 130 213 188 225
rect 288 331 346 343
rect 288 225 300 331
rect 334 225 346 331
rect 288 213 346 225
<< mvpdiff >>
rect 130 1821 188 1833
rect 130 1645 142 1821
rect 176 1645 188 1821
rect 130 1633 188 1645
rect 288 1821 346 1833
rect 288 1645 300 1821
rect 334 1645 346 1821
rect 288 1633 346 1645
rect 130 1385 188 1397
rect 130 1209 142 1385
rect 176 1209 188 1385
rect 130 1197 188 1209
rect 288 1385 346 1397
rect 288 1209 300 1385
rect 334 1209 346 1385
rect 288 1197 346 1209
<< mvndiffc >>
rect 142 573 176 679
rect 300 573 334 679
rect 142 225 176 331
rect 300 225 334 331
<< mvpdiffc >>
rect 142 1645 176 1821
rect 300 1645 334 1821
rect 142 1209 176 1385
rect 300 1209 334 1385
<< mvpsubdiff >>
rect -2 856 488 868
rect -2 822 124 856
rect 352 822 488 856
rect -2 810 488 822
rect -2 760 56 810
rect -2 144 10 760
rect 44 144 56 760
rect 430 760 488 810
rect -2 94 56 144
rect 430 144 442 760
rect 476 144 488 760
rect 430 94 488 144
rect -2 82 488 94
rect -2 48 124 82
rect 352 48 488 82
rect -2 36 488 48
<< mvnsubdiff >>
rect 18 1998 458 2010
rect 18 1964 124 1998
rect 352 1964 458 1998
rect 18 1952 458 1964
rect 18 1902 76 1952
rect 18 1128 30 1902
rect 64 1128 76 1902
rect 400 1902 458 1952
rect 18 1078 76 1128
rect 400 1128 412 1902
rect 446 1128 458 1902
rect 400 1078 458 1128
rect 18 1066 458 1078
rect 18 1032 124 1066
rect 352 1032 458 1066
rect 18 1020 458 1032
<< mvpsubdiffcont >>
rect 124 822 352 856
rect 10 144 44 760
rect 442 144 476 760
rect 124 48 352 82
<< mvnsubdiffcont >>
rect 124 1964 352 1998
rect 30 1128 64 1902
rect 412 1128 446 1902
rect 124 1032 352 1066
<< poly >>
rect 188 1914 288 1930
rect 188 1880 204 1914
rect 272 1880 288 1914
rect 188 1833 288 1880
rect 188 1586 288 1633
rect 188 1552 204 1586
rect 272 1552 288 1586
rect 188 1536 288 1552
rect 188 1478 288 1494
rect 188 1444 204 1478
rect 272 1444 288 1478
rect 188 1397 288 1444
rect 188 1150 288 1197
rect 188 1116 204 1150
rect 272 1116 288 1150
rect 188 1100 288 1116
rect 188 763 288 779
rect 188 729 204 763
rect 272 729 288 763
rect 188 691 288 729
rect 188 523 288 561
rect 188 489 204 523
rect 272 489 288 523
rect 188 473 288 489
rect 188 415 288 431
rect 188 381 204 415
rect 272 381 288 415
rect 188 343 288 381
rect 188 175 288 213
rect 188 141 204 175
rect 272 141 288 175
rect 188 125 288 141
<< polycont >>
rect 204 1880 272 1914
rect 204 1552 272 1586
rect 204 1444 272 1478
rect 204 1116 272 1150
rect 204 729 272 763
rect 204 489 272 523
rect 204 381 272 415
rect 204 141 272 175
<< locali >>
rect 30 1964 124 1998
rect 352 1964 446 1998
rect 30 1902 64 1964
rect 188 1880 204 1914
rect 272 1880 288 1914
rect 412 1902 446 1964
rect 142 1821 176 1837
rect 142 1629 176 1645
rect 300 1821 334 1837
rect 300 1629 334 1645
rect 188 1552 204 1586
rect 272 1552 288 1586
rect 188 1444 204 1478
rect 272 1444 288 1478
rect 142 1385 176 1401
rect 142 1193 176 1209
rect 300 1385 334 1401
rect 300 1193 334 1209
rect 30 1066 64 1128
rect 188 1116 204 1150
rect 272 1116 288 1150
rect 412 1066 446 1128
rect 30 1032 124 1066
rect 352 1032 446 1066
rect 10 822 124 856
rect 352 822 476 856
rect 10 760 44 822
rect 188 729 204 763
rect 272 729 288 763
rect 442 760 476 822
rect 142 679 176 695
rect 142 557 176 573
rect 300 679 334 695
rect 300 557 334 573
rect 188 489 204 523
rect 272 489 288 523
rect 188 381 204 415
rect 272 381 288 415
rect 142 331 176 347
rect 142 209 176 225
rect 300 331 334 347
rect 300 209 334 225
rect 10 82 44 144
rect 188 141 204 175
rect 272 141 288 175
rect 442 82 476 144
rect 10 48 124 82
rect 352 48 476 82
<< viali >>
rect 124 1964 352 1998
rect 204 1880 272 1914
rect 142 1645 176 1821
rect 300 1645 334 1821
rect 204 1552 272 1586
rect 204 1444 272 1478
rect 142 1209 176 1385
rect 300 1209 334 1385
rect 204 1116 272 1150
rect 204 729 272 763
rect 142 573 176 679
rect 300 573 334 679
rect 204 489 272 523
rect 204 381 272 415
rect 142 225 176 331
rect 300 225 334 331
rect 204 141 272 175
rect 124 48 352 82
<< metal1 >>
rect 100 1998 376 2010
rect 100 1964 124 1998
rect 352 1964 376 1998
rect 100 1952 376 1964
rect 192 1914 284 1920
rect 192 1880 204 1914
rect 272 1880 284 1914
rect 192 1874 284 1880
rect 136 1821 182 1833
rect 136 1645 142 1821
rect 176 1645 182 1821
rect 136 1633 182 1645
rect 221 1592 255 1874
rect 294 1821 340 1833
rect 294 1645 300 1821
rect 334 1645 340 1821
rect 294 1633 340 1645
rect 192 1586 284 1592
rect 192 1552 204 1586
rect 272 1552 284 1586
rect 192 1546 284 1552
rect 192 1478 284 1484
rect 192 1444 204 1478
rect 272 1444 284 1478
rect 192 1438 284 1444
rect 136 1385 182 1397
rect 136 1209 142 1385
rect 176 1209 182 1385
rect 136 1197 182 1209
rect 221 1156 255 1438
rect 294 1385 340 1397
rect 294 1209 300 1385
rect 334 1209 340 1385
rect 294 1197 340 1209
rect 192 1150 284 1156
rect 192 1116 204 1150
rect 272 1116 284 1150
rect 192 1110 284 1116
rect 192 763 284 769
rect 192 729 204 763
rect 272 729 284 763
rect 192 723 284 729
rect 136 679 182 691
rect 136 573 142 679
rect 176 573 182 679
rect 136 561 182 573
rect 221 529 255 723
rect 294 679 340 691
rect 294 573 300 679
rect 334 573 340 679
rect 294 561 340 573
rect 192 523 284 529
rect 192 489 204 523
rect 272 489 284 523
rect 192 483 284 489
rect 192 415 284 421
rect 192 381 204 415
rect 272 381 284 415
rect 192 375 284 381
rect 136 331 182 343
rect 136 225 142 331
rect 176 225 182 331
rect 136 213 182 225
rect 221 181 255 375
rect 294 331 340 343
rect 294 225 300 331
rect 334 225 340 331
rect 294 213 340 225
rect 192 175 284 181
rect 192 141 204 175
rect 272 141 284 175
rect 192 135 284 141
rect 100 82 376 94
rect 100 48 124 82
rect 352 48 376 82
rect 100 36 376 48
<< labels >>
flabel metal1 100 1952 376 2010 0 FreeSans 256 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal1 100 36 376 94 0 FreeSans 256 0 0 0 VSS
port 2 nsew ground bidirectional
<< end >>
