magic
tech sky130A
magscale 1 2
timestamp 1727607685
<< metal1 >>
rect 88 6003 388 6061
rect 221 5019 255 5971
rect 297 5051 303 5103
rect 355 5051 361 5103
rect 206 4967 212 5019
rect 264 4967 270 5019
rect 88 4871 388 4929
rect 88 2510 388 2568
rect 130 2187 164 2510
rect 212 2095 264 2159
rect 121 2031 173 2037
rect 121 1973 173 1979
rect 130 1757 164 1973
rect 221 1847 255 2095
rect 206 1795 212 1847
rect 264 1795 270 1847
rect 130 1723 254 1757
rect 130 1436 164 1689
rect 312 1616 346 2395
rect 303 1610 355 1616
rect 303 1552 355 1558
rect 312 1551 346 1552
rect 88 1378 388 1436
rect 88 1168 388 1226
rect 130 845 164 1168
rect 316 1130 322 1139
rect 220 1096 322 1130
rect 316 1087 322 1096
rect 374 1087 380 1139
rect 312 1042 346 1053
rect 297 990 303 1042
rect 355 990 361 1042
rect 212 424 264 430
rect 212 366 264 372
rect 130 94 164 347
rect 312 209 346 990
rect 88 36 388 94
<< via1 >>
rect 303 5051 355 5103
rect 212 4967 264 5019
rect 121 1979 173 2031
rect 212 1795 264 1847
rect 303 1558 355 1610
rect 322 1087 374 1139
rect 303 990 355 1042
rect 212 372 264 424
<< metal2 >>
rect 303 5103 355 5109
rect 303 5045 355 5051
rect 212 5019 264 5025
rect 212 4961 264 4967
rect 115 1979 121 2031
rect 173 2022 179 2031
rect 221 2022 255 4961
rect 173 1988 255 2022
rect 173 1979 179 1988
rect 312 1929 346 5045
rect 130 1895 346 1929
rect 130 595 164 1895
rect 212 1847 264 1853
rect 212 1789 264 1795
rect 221 1033 255 1789
rect 297 1558 303 1610
rect 355 1558 361 1610
rect 312 1145 346 1558
rect 312 1139 374 1145
rect 312 1096 322 1139
rect 322 1081 374 1087
rect 303 1042 355 1048
rect 221 999 303 1033
rect 303 984 355 990
rect 130 561 255 595
rect 221 424 255 561
rect 206 372 212 424
rect 264 372 270 424
use inverter  inverter_0
timestamp 1727607685
transform 1 0 0 0 1 4835
box 0 0 476 1292
use transistor_pair  transistor_pair_0
timestamp 1727597281
transform 1 0 0 0 1 1342
box 0 0 476 1292
use transistor_pair  transistor_pair_1
timestamp 1727597281
transform 1 0 0 0 1 0
box 0 0 476 1292
<< labels >>
flabel metal1 312 209 346 1053 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 88 2510 388 2568 0 FreeSans 256 0 0 0 OVDD1
port 3 nsew
flabel metal1 88 1378 388 1436 0 FreeSans 256 0 0 0 VSS1
port 6 nsew
flabel metal1 88 1168 388 1226 0 FreeSans 256 0 0 0 OVDD2
port 4 nsew
flabel metal1 88 36 388 94 0 FreeSans 256 0 0 0 VSS2
port 7 nsew
flabel metal1 221 4976 255 5965 0 FreeSans 256 0 0 0 IN
port 0 nsew
flabel metal1 88 4871 388 4929 0 FreeSans 256 0 0 0 VSS0
port 5 nsew
flabel metal1 88 6003 388 6061 0 FreeSans 256 0 0 0 IVDD
port 1 nsew
<< end >>
