magic
tech sky130A
magscale 1 2
timestamp 1731100676
<< dnwell >>
rect -301 -335 3907 13976
<< nwell >>
rect -381 13770 3987 14056
rect -381 -129 -95 13770
rect 3701 -129 3987 13770
rect -381 -415 3987 -129
<< nsubdiff >>
rect -344 13999 3950 14019
rect -344 13965 -264 13999
rect 3870 13965 3950 13999
rect -344 13945 3950 13965
rect -344 13939 -270 13945
rect -344 -298 -324 13939
rect -290 -298 -270 13939
rect -344 -304 -270 -298
rect 3876 13939 3950 13945
rect 3876 -298 3896 13939
rect 3930 -298 3950 13939
rect 3876 -304 3950 -298
rect -344 -324 3950 -304
rect -344 -358 -264 -324
rect 3870 -358 3950 -324
rect -344 -378 3950 -358
<< nsubdiffcont >>
rect -264 13965 3870 13999
rect -324 -298 -290 13939
rect 3896 -298 3930 13939
rect -264 -358 3870 -324
<< locali >>
rect -324 13965 -264 13999
rect 3870 13965 3930 13999
rect -324 13939 -290 13965
rect -324 -324 -290 -298
rect 3896 13939 3930 13965
rect 3896 -324 3930 -298
rect -324 -358 -264 -324
rect 3870 -358 3930 -324
use decoder4_signed  decoder4_signed_0
timestamp 1731100676
transform 1 0 305 0 1 0
box -305 0 2996 13410
<< end >>
