magic
tech sky130A
magscale 1 2
timestamp 1727605625
<< dnwell >>
rect -654 -335 1130 2682
<< nwell >>
rect -734 2476 1210 2762
rect -734 -129 -448 2476
rect 924 -129 1210 2476
rect -734 -415 1210 -129
<< nsubdiff >>
rect -697 2705 1173 2725
rect -697 2671 -617 2705
rect 1093 2671 1173 2705
rect -697 2651 1173 2671
rect -697 2645 -623 2651
rect -697 -298 -677 2645
rect -643 -298 -623 2645
rect -697 -304 -623 -298
rect 1099 2645 1173 2651
rect 1099 -298 1119 2645
rect 1153 -298 1173 2645
rect 1099 -304 1173 -298
rect -697 -324 1173 -304
rect -697 -358 -617 -324
rect 1093 -358 1173 -324
rect -697 -378 1173 -358
<< nsubdiffcont >>
rect -617 2671 1093 2705
rect -677 -298 -643 2645
rect 1119 -298 1153 2645
rect -617 -358 1093 -324
<< locali >>
rect -677 2671 -617 2705
rect 1093 2671 1153 2705
rect -677 2645 -643 2671
rect -677 -324 -643 -298
rect 1119 2645 1153 2671
rect 1119 -324 1153 -298
rect -677 -358 -617 -324
rect 1093 -358 1153 -324
use passgate_single  passgate_single_0
timestamp 1727605497
transform 1 0 0 0 1 0
box -48 0 524 2076
<< end >>
