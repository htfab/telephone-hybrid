magic
tech sky130A
timestamp 1727641773
use tie_high  tie_high_1
array 0 7 150 0 0 646
timestamp 1727638007
transform 1 0 0 0 1 0
box 44 18 194 613
use transistor_pair_bus  transistor_pair_bus_0
timestamp 1727637843
transform 1 0 0 0 1 0
box -30 0 1318 646
<< end >>
