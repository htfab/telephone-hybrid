magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< xpolycontact >>
rect -2110 3184 -2040 3616
rect -2110 -3616 -2040 -3184
rect -1944 3184 -1874 3616
rect -1944 -3616 -1874 -3184
rect -1778 3184 -1708 3616
rect -1778 -3616 -1708 -3184
rect -1612 3184 -1542 3616
rect -1612 -3616 -1542 -3184
rect -1446 3184 -1376 3616
rect -1446 -3616 -1376 -3184
rect -1280 3184 -1210 3616
rect -1280 -3616 -1210 -3184
rect -1114 3184 -1044 3616
rect -1114 -3616 -1044 -3184
rect -948 3184 -878 3616
rect -948 -3616 -878 -3184
rect -782 3184 -712 3616
rect -782 -3616 -712 -3184
rect -616 3184 -546 3616
rect -616 -3616 -546 -3184
rect -450 3184 -380 3616
rect -450 -3616 -380 -3184
rect -284 3184 -214 3616
rect -284 -3616 -214 -3184
rect -118 3184 -48 3616
rect -118 -3616 -48 -3184
rect 48 3184 118 3616
rect 48 -3616 118 -3184
rect 214 3184 284 3616
rect 214 -3616 284 -3184
rect 380 3184 450 3616
rect 380 -3616 450 -3184
rect 546 3184 616 3616
rect 546 -3616 616 -3184
rect 712 3184 782 3616
rect 712 -3616 782 -3184
rect 878 3184 948 3616
rect 878 -3616 948 -3184
rect 1044 3184 1114 3616
rect 1044 -3616 1114 -3184
rect 1210 3184 1280 3616
rect 1210 -3616 1280 -3184
rect 1376 3184 1446 3616
rect 1376 -3616 1446 -3184
rect 1542 3184 1612 3616
rect 1542 -3616 1612 -3184
rect 1708 3184 1778 3616
rect 1708 -3616 1778 -3184
rect 1874 3184 1944 3616
rect 1874 -3616 1944 -3184
rect 2040 3184 2110 3616
rect 2040 -3616 2110 -3184
<< xpolyres >>
rect -2110 -3184 -2040 3184
rect -1944 -3184 -1874 3184
rect -1778 -3184 -1708 3184
rect -1612 -3184 -1542 3184
rect -1446 -3184 -1376 3184
rect -1280 -3184 -1210 3184
rect -1114 -3184 -1044 3184
rect -948 -3184 -878 3184
rect -782 -3184 -712 3184
rect -616 -3184 -546 3184
rect -450 -3184 -380 3184
rect -284 -3184 -214 3184
rect -118 -3184 -48 3184
rect 48 -3184 118 3184
rect 214 -3184 284 3184
rect 380 -3184 450 3184
rect 546 -3184 616 3184
rect 712 -3184 782 3184
rect 878 -3184 948 3184
rect 1044 -3184 1114 3184
rect 1210 -3184 1280 3184
rect 1376 -3184 1446 3184
rect 1542 -3184 1612 3184
rect 1708 -3184 1778 3184
rect 1874 -3184 1944 3184
rect 2040 -3184 2110 3184
<< viali >>
rect -2094 3201 -2056 3598
rect -1928 3201 -1890 3598
rect -1762 3201 -1724 3598
rect -1596 3201 -1558 3598
rect -1430 3201 -1392 3598
rect -1264 3201 -1226 3598
rect -1098 3201 -1060 3598
rect -932 3201 -894 3598
rect -766 3201 -728 3598
rect -600 3201 -562 3598
rect -434 3201 -396 3598
rect -268 3201 -230 3598
rect -102 3201 -64 3598
rect 64 3201 102 3598
rect 230 3201 268 3598
rect 396 3201 434 3598
rect 562 3201 600 3598
rect 728 3201 766 3598
rect 894 3201 932 3598
rect 1060 3201 1098 3598
rect 1226 3201 1264 3598
rect 1392 3201 1430 3598
rect 1558 3201 1596 3598
rect 1724 3201 1762 3598
rect 1890 3201 1928 3598
rect 2056 3201 2094 3598
rect -2094 -3598 -2056 -3201
rect -1928 -3598 -1890 -3201
rect -1762 -3598 -1724 -3201
rect -1596 -3598 -1558 -3201
rect -1430 -3598 -1392 -3201
rect -1264 -3598 -1226 -3201
rect -1098 -3598 -1060 -3201
rect -932 -3598 -894 -3201
rect -766 -3598 -728 -3201
rect -600 -3598 -562 -3201
rect -434 -3598 -396 -3201
rect -268 -3598 -230 -3201
rect -102 -3598 -64 -3201
rect 64 -3598 102 -3201
rect 230 -3598 268 -3201
rect 396 -3598 434 -3201
rect 562 -3598 600 -3201
rect 728 -3598 766 -3201
rect 894 -3598 932 -3201
rect 1060 -3598 1098 -3201
rect 1226 -3598 1264 -3201
rect 1392 -3598 1430 -3201
rect 1558 -3598 1596 -3201
rect 1724 -3598 1762 -3201
rect 1890 -3598 1928 -3201
rect 2056 -3598 2094 -3201
<< metal1 >>
rect -2100 3598 -2050 3610
rect -2100 3201 -2094 3598
rect -2056 3201 -2050 3598
rect -2100 3189 -2050 3201
rect -1934 3598 -1884 3610
rect -1934 3201 -1928 3598
rect -1890 3201 -1884 3598
rect -1934 3189 -1884 3201
rect -1768 3598 -1718 3610
rect -1768 3201 -1762 3598
rect -1724 3201 -1718 3598
rect -1768 3189 -1718 3201
rect -1602 3598 -1552 3610
rect -1602 3201 -1596 3598
rect -1558 3201 -1552 3598
rect -1602 3189 -1552 3201
rect -1436 3598 -1386 3610
rect -1436 3201 -1430 3598
rect -1392 3201 -1386 3598
rect -1436 3189 -1386 3201
rect -1270 3598 -1220 3610
rect -1270 3201 -1264 3598
rect -1226 3201 -1220 3598
rect -1270 3189 -1220 3201
rect -1104 3598 -1054 3610
rect -1104 3201 -1098 3598
rect -1060 3201 -1054 3598
rect -1104 3189 -1054 3201
rect -938 3598 -888 3610
rect -938 3201 -932 3598
rect -894 3201 -888 3598
rect -938 3189 -888 3201
rect -772 3598 -722 3610
rect -772 3201 -766 3598
rect -728 3201 -722 3598
rect -772 3189 -722 3201
rect -606 3598 -556 3610
rect -606 3201 -600 3598
rect -562 3201 -556 3598
rect -606 3189 -556 3201
rect -440 3598 -390 3610
rect -440 3201 -434 3598
rect -396 3201 -390 3598
rect -440 3189 -390 3201
rect -274 3598 -224 3610
rect -274 3201 -268 3598
rect -230 3201 -224 3598
rect -274 3189 -224 3201
rect -108 3598 -58 3610
rect -108 3201 -102 3598
rect -64 3201 -58 3598
rect -108 3189 -58 3201
rect 58 3598 108 3610
rect 58 3201 64 3598
rect 102 3201 108 3598
rect 58 3189 108 3201
rect 224 3598 274 3610
rect 224 3201 230 3598
rect 268 3201 274 3598
rect 224 3189 274 3201
rect 390 3598 440 3610
rect 390 3201 396 3598
rect 434 3201 440 3598
rect 390 3189 440 3201
rect 556 3598 606 3610
rect 556 3201 562 3598
rect 600 3201 606 3598
rect 556 3189 606 3201
rect 722 3598 772 3610
rect 722 3201 728 3598
rect 766 3201 772 3598
rect 722 3189 772 3201
rect 888 3598 938 3610
rect 888 3201 894 3598
rect 932 3201 938 3598
rect 888 3189 938 3201
rect 1054 3598 1104 3610
rect 1054 3201 1060 3598
rect 1098 3201 1104 3598
rect 1054 3189 1104 3201
rect 1220 3598 1270 3610
rect 1220 3201 1226 3598
rect 1264 3201 1270 3598
rect 1220 3189 1270 3201
rect 1386 3598 1436 3610
rect 1386 3201 1392 3598
rect 1430 3201 1436 3598
rect 1386 3189 1436 3201
rect 1552 3598 1602 3610
rect 1552 3201 1558 3598
rect 1596 3201 1602 3598
rect 1552 3189 1602 3201
rect 1718 3598 1768 3610
rect 1718 3201 1724 3598
rect 1762 3201 1768 3598
rect 1718 3189 1768 3201
rect 1884 3598 1934 3610
rect 1884 3201 1890 3598
rect 1928 3201 1934 3598
rect 1884 3189 1934 3201
rect 2050 3598 2100 3610
rect 2050 3201 2056 3598
rect 2094 3201 2100 3598
rect 2050 3189 2100 3201
rect -2100 -3201 -2050 -3189
rect -2100 -3598 -2094 -3201
rect -2056 -3598 -2050 -3201
rect -2100 -3610 -2050 -3598
rect -1934 -3201 -1884 -3189
rect -1934 -3598 -1928 -3201
rect -1890 -3598 -1884 -3201
rect -1934 -3610 -1884 -3598
rect -1768 -3201 -1718 -3189
rect -1768 -3598 -1762 -3201
rect -1724 -3598 -1718 -3201
rect -1768 -3610 -1718 -3598
rect -1602 -3201 -1552 -3189
rect -1602 -3598 -1596 -3201
rect -1558 -3598 -1552 -3201
rect -1602 -3610 -1552 -3598
rect -1436 -3201 -1386 -3189
rect -1436 -3598 -1430 -3201
rect -1392 -3598 -1386 -3201
rect -1436 -3610 -1386 -3598
rect -1270 -3201 -1220 -3189
rect -1270 -3598 -1264 -3201
rect -1226 -3598 -1220 -3201
rect -1270 -3610 -1220 -3598
rect -1104 -3201 -1054 -3189
rect -1104 -3598 -1098 -3201
rect -1060 -3598 -1054 -3201
rect -1104 -3610 -1054 -3598
rect -938 -3201 -888 -3189
rect -938 -3598 -932 -3201
rect -894 -3598 -888 -3201
rect -938 -3610 -888 -3598
rect -772 -3201 -722 -3189
rect -772 -3598 -766 -3201
rect -728 -3598 -722 -3201
rect -772 -3610 -722 -3598
rect -606 -3201 -556 -3189
rect -606 -3598 -600 -3201
rect -562 -3598 -556 -3201
rect -606 -3610 -556 -3598
rect -440 -3201 -390 -3189
rect -440 -3598 -434 -3201
rect -396 -3598 -390 -3201
rect -440 -3610 -390 -3598
rect -274 -3201 -224 -3189
rect -274 -3598 -268 -3201
rect -230 -3598 -224 -3201
rect -274 -3610 -224 -3598
rect -108 -3201 -58 -3189
rect -108 -3598 -102 -3201
rect -64 -3598 -58 -3201
rect -108 -3610 -58 -3598
rect 58 -3201 108 -3189
rect 58 -3598 64 -3201
rect 102 -3598 108 -3201
rect 58 -3610 108 -3598
rect 224 -3201 274 -3189
rect 224 -3598 230 -3201
rect 268 -3598 274 -3201
rect 224 -3610 274 -3598
rect 390 -3201 440 -3189
rect 390 -3598 396 -3201
rect 434 -3598 440 -3201
rect 390 -3610 440 -3598
rect 556 -3201 606 -3189
rect 556 -3598 562 -3201
rect 600 -3598 606 -3201
rect 556 -3610 606 -3598
rect 722 -3201 772 -3189
rect 722 -3598 728 -3201
rect 766 -3598 772 -3201
rect 722 -3610 772 -3598
rect 888 -3201 938 -3189
rect 888 -3598 894 -3201
rect 932 -3598 938 -3201
rect 888 -3610 938 -3598
rect 1054 -3201 1104 -3189
rect 1054 -3598 1060 -3201
rect 1098 -3598 1104 -3201
rect 1054 -3610 1104 -3598
rect 1220 -3201 1270 -3189
rect 1220 -3598 1226 -3201
rect 1264 -3598 1270 -3201
rect 1220 -3610 1270 -3598
rect 1386 -3201 1436 -3189
rect 1386 -3598 1392 -3201
rect 1430 -3598 1436 -3201
rect 1386 -3610 1436 -3598
rect 1552 -3201 1602 -3189
rect 1552 -3598 1558 -3201
rect 1596 -3598 1602 -3201
rect 1552 -3610 1602 -3598
rect 1718 -3201 1768 -3189
rect 1718 -3598 1724 -3201
rect 1762 -3598 1768 -3201
rect 1718 -3610 1768 -3598
rect 1884 -3201 1934 -3189
rect 1884 -3598 1890 -3201
rect 1928 -3598 1934 -3201
rect 1884 -3610 1934 -3598
rect 2050 -3201 2100 -3189
rect 2050 -3598 2056 -3201
rect 2094 -3598 2100 -3201
rect 2050 -3610 2100 -3598
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 32.0 m 1 nx 26 wmin 0.350 lmin 0.50 rho 2000 val 183.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
