magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< metal1 >>
rect 3204 6959 3440 7391
rect 3536 6959 3772 7391
rect 3868 6959 4104 7391
rect 4200 6959 4436 7391
rect 4532 6959 4768 7391
rect 4864 6959 5100 7391
rect 5196 6959 5432 7391
rect 5528 6959 5764 7391
rect 5860 6959 6096 7391
rect 6192 6959 6428 7391
rect 6524 6959 6760 7391
rect 6856 6959 7092 7391
rect 3204 574 3274 591
rect 3204 177 3213 574
rect 3265 177 3274 574
rect 3204 159 3274 177
rect 3370 159 3606 591
rect 3702 159 3938 591
rect 4034 159 4270 591
rect 4366 463 4602 591
rect 4366 287 4390 463
rect 4578 287 4602 463
rect 4366 159 4602 287
rect 4698 159 4934 591
rect 5030 159 5266 591
rect 5362 159 5598 591
rect 5694 463 5930 591
rect 5694 287 5718 463
rect 5906 287 5930 463
rect 5694 159 5930 287
rect 6026 159 6262 591
rect 6358 159 6594 591
rect 6690 159 6926 591
rect 7022 574 7092 591
rect 7022 177 7031 574
rect 7083 177 7092 574
rect 7022 159 7092 177
rect 5434 -6 5626 0
rect 5434 -58 5446 -6
rect 5614 -58 5626 -6
rect 5434 -64 5626 -58
rect 5810 -6 6002 0
rect 5810 -58 5822 -6
rect 5990 -58 6002 -6
rect 5810 -64 6002 -58
<< via1 >>
rect 3213 177 3265 574
rect 4390 287 4578 463
rect 5718 287 5906 463
rect 7031 177 7083 574
rect 5446 -58 5614 -6
rect 5822 -58 5990 -6
<< metal2 >>
rect 3204 574 3274 591
rect 3204 177 3213 574
rect 3265 177 3274 574
rect 7022 574 7092 591
rect 4384 463 4584 475
rect 4384 287 4390 463
rect 4578 287 4584 463
rect 4384 275 4584 287
rect 5706 463 5918 469
rect 5706 287 5718 463
rect 5906 287 5918 463
rect 5706 281 5918 287
rect 3204 159 3274 177
rect 3215 120 3263 159
rect 5787 120 5836 281
rect 7022 177 7031 574
rect 7083 177 7092 574
rect 7022 159 7092 177
rect 7032 120 7080 159
rect 3215 72 5554 120
rect 5506 0 5554 72
rect 5787 71 5931 120
rect 6084 72 7080 120
rect 5882 0 5930 71
rect 5434 -6 5626 0
rect 5434 -58 5446 -6
rect 5614 -58 5626 -6
rect 5434 -64 5626 -58
rect 5810 -6 6002 0
rect 5810 -58 5822 -6
rect 5990 -58 6002 -6
rect 5810 -64 6002 -58
rect 6084 -1930 6132 72
rect 3204 -2248 3404 -2048
rect 3204 -2506 3404 -2306
rect 3204 -3022 3404 -2822
rect 3204 -3276 3404 -3076
use sky130_fd_pr__res_xhigh_po_0p35_H47ZCG  sky130_fd_pr__res_xhigh_po_0p35_H47ZCG_0
timestamp 1727597281
transform 1 0 6476 0 1 3775
box -616 -3616 616 3616
use opamp  x1
timestamp 1727597281
transform 1 0 0 0 1 -1600
box 3204 -1676 6132 1720
use sky130_fd_pr__res_xhigh_po_0p35_H47ZCG  XR1
timestamp 1727597281
transform 1 0 3820 0 1 3775
box -616 -3616 616 3616
use sky130_fd_pr__res_xhigh_po_0p35_H47ZCG  XR2
timestamp 1727597281
transform 1 0 5148 0 1 3775
box -616 -3616 616 3616
<< labels >>
flabel metal2 3204 -3022 3404 -2822 0 FreeSans 128 0 0 0 OUT
port 2 nsew
flabel metal2 3204 -3276 3404 -3076 0 FreeSans 128 0 0 0 VSS
port 4 nsew
flabel metal2 3204 -2248 3404 -2048 0 FreeSans 128 0 0 0 VDD
port 3 nsew
flabel metal2 3204 -2506 3404 -2306 0 FreeSans 128 0 0 0 LINE
port 1 nsew
flabel metal2 4384 275 4584 475 0 FreeSans 128 0 0 0 IN
port 0 nsew
<< end >>
