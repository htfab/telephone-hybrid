magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< nwell >>
rect 0 606 476 1292
<< pwell >>
rect 0 0 476 556
<< mvpsubdiff >>
rect 88 508 388 520
rect 88 474 124 508
rect 352 474 388 508
rect 88 462 388 474
rect 88 82 388 94
rect 88 48 124 82
rect 352 48 388 82
rect 88 36 388 48
<< mvnsubdiff >>
rect 88 1214 388 1226
rect 88 1180 124 1214
rect 352 1180 388 1214
rect 88 1168 388 1180
rect 88 718 388 730
rect 88 684 124 718
rect 352 684 388 718
rect 88 672 388 684
<< mvpsubdiffcont >>
rect 124 474 352 508
rect 124 48 352 82
<< mvnsubdiffcont >>
rect 124 1180 352 1214
rect 124 684 352 718
<< locali >>
rect 88 1180 124 1214
rect 352 1180 388 1214
rect 88 684 124 718
rect 352 684 388 718
rect 88 474 124 508
rect 352 474 388 508
rect 88 48 124 82
rect 352 48 388 82
<< viali >>
rect 124 1180 352 1214
rect 124 48 352 82
<< metal1 >>
rect 88 1214 388 1226
rect 88 1180 124 1214
rect 352 1180 388 1214
rect 88 1168 388 1180
rect 130 845 164 1053
rect 221 768 255 1130
rect 312 845 346 1053
rect 130 209 164 347
rect 221 141 255 415
rect 312 209 346 347
rect 88 82 388 94
rect 88 48 124 82
rect 352 48 388 82
rect 88 36 388 48
use nfet  nfet_0
timestamp 1727597281
transform 1 0 238 0 1 278
box -120 -153 120 153
use pfet  pfet_0
timestamp 1727597281
transform 1 0 238 0 1 949
box -186 -200 186 200
<< end >>
