magic
tech sky130A
magscale 1 2
timestamp 1731100676
<< metal1 >>
rect 203 2509 209 2569
rect 269 2509 275 2569
rect 803 2509 809 2569
rect 869 2509 875 2569
rect 1403 2509 1409 2569
rect 1469 2509 1475 2569
rect 2003 2509 2009 2569
rect 2069 2509 2075 2569
rect 2603 2509 2609 2569
rect 2669 2509 2675 2569
rect 1766 2343 1772 2395
rect 1824 2343 1830 2395
rect 2666 2343 2672 2395
rect 2724 2343 2730 2395
rect 1466 2259 1472 2311
rect 1524 2259 1530 2311
rect 2366 2175 2372 2227
rect 2424 2175 2430 2227
rect 2366 2150 2430 2175
rect 738 2133 744 2142
rect 672 2099 744 2133
rect 738 2090 744 2099
rect 796 2090 802 2142
rect 1166 2091 1172 2143
rect 1224 2091 1230 2143
rect 2066 2091 2072 2143
rect 2124 2091 2130 2143
rect 572 1964 624 1970
rect 657 1912 663 1964
rect 715 1912 721 1964
rect 866 1912 872 1964
rect 924 1912 930 1964
rect 572 1906 624 1912
rect 957 1551 963 1603
rect 1015 1551 1021 1603
rect 281 1507 314 1511
rect 281 1390 315 1507
rect 503 1377 509 1437
rect 569 1377 575 1437
rect 1103 1377 1109 1437
rect 1169 1377 1175 1437
rect 1703 1377 1709 1437
rect 1769 1377 1775 1437
rect 2303 1377 2309 1437
rect 2369 1377 2375 1437
rect 203 1167 209 1227
rect 269 1167 275 1227
rect 803 1167 809 1227
rect 869 1167 875 1227
rect 1403 1167 1409 1227
rect 1469 1167 1475 1227
rect 2003 1167 2009 1227
rect 2069 1167 2075 1227
rect 2603 1167 2609 1227
rect 2669 1167 2675 1227
rect 357 1001 363 1053
rect 415 1001 421 1053
rect 1766 1001 1772 1053
rect 1824 1001 1830 1053
rect 2666 1001 2672 1053
rect 2724 1001 2730 1053
rect 957 917 963 969
rect 1015 917 1021 969
rect 1466 917 1472 969
rect 1524 917 1530 969
rect 657 833 663 885
rect 715 833 721 885
rect 2366 833 2372 885
rect 2424 833 2430 885
rect 2366 808 2430 833
rect 1166 749 1172 801
rect 1224 749 1230 801
rect 2066 749 2072 801
rect 2124 749 2130 801
rect 572 622 624 628
rect 657 570 663 622
rect 715 570 721 622
rect 866 570 872 622
rect 924 570 930 622
rect 572 564 624 570
rect 266 209 272 261
rect 324 209 330 261
rect 503 35 509 95
rect 569 35 575 95
rect 1103 35 1109 95
rect 1169 35 1175 95
rect 1703 35 1709 95
rect 1769 35 1775 95
rect 2303 35 2309 95
rect 2369 35 2375 95
<< via1 >>
rect 209 2509 269 2569
rect 809 2509 869 2569
rect 1409 2509 1469 2569
rect 2009 2509 2069 2569
rect 2609 2509 2669 2569
rect 1772 2343 1824 2395
rect 2672 2343 2724 2395
rect 1472 2259 1524 2311
rect 2372 2175 2424 2227
rect 744 2090 796 2142
rect 1172 2091 1224 2143
rect 2072 2091 2124 2143
rect 572 1912 624 1964
rect 663 1912 715 1964
rect 872 1912 924 1964
rect 963 1551 1015 1603
rect 509 1377 569 1437
rect 1109 1377 1169 1437
rect 1709 1377 1769 1437
rect 2309 1377 2369 1437
rect 209 1167 269 1227
rect 809 1167 869 1227
rect 1409 1167 1469 1227
rect 2009 1167 2069 1227
rect 2609 1167 2669 1227
rect 363 1001 415 1053
rect 1772 1001 1824 1053
rect 2672 1001 2724 1053
rect 963 917 1015 969
rect 1472 917 1524 969
rect 663 833 715 885
rect 2372 833 2424 885
rect 1172 749 1224 801
rect 2072 749 2124 801
rect 572 570 624 622
rect 663 570 715 622
rect 872 570 924 622
rect 272 209 324 261
rect 509 35 569 95
rect 1109 35 1169 95
rect 1709 35 1769 95
rect 2309 35 2369 95
<< metal2 >>
rect 209 2569 269 2578
rect 209 2500 269 2509
rect 809 2569 869 2578
rect 809 2500 869 2509
rect 1409 2569 1469 2578
rect 1409 2500 1469 2509
rect 2009 2569 2069 2578
rect 2009 2500 2069 2509
rect 2609 2569 2669 2578
rect 2609 2500 2669 2509
rect 359 2399 419 2408
rect 1772 2395 1824 2401
rect 419 2352 1772 2386
rect 359 2330 419 2339
rect 2672 2395 2724 2401
rect 1824 2352 2672 2386
rect 1772 2337 1824 2343
rect 2672 2337 2724 2343
rect 959 2315 1019 2324
rect 1472 2311 1524 2317
rect 1019 2268 1472 2302
rect 959 2246 1019 2255
rect 1472 2253 1524 2259
rect 659 2231 719 2240
rect 2372 2227 2424 2233
rect 719 2184 2372 2218
rect 659 2162 719 2171
rect 2372 2169 2424 2175
rect 744 2142 796 2148
rect 672 2100 744 2134
rect 1172 2143 1224 2149
rect 796 2100 1172 2134
rect 744 2084 796 2090
rect 2072 2143 2124 2149
rect 1224 2100 2072 2134
rect 1172 2085 1224 2091
rect 2072 2085 2124 2091
rect 663 1964 715 1970
rect 566 1955 572 1964
rect 148 1921 572 1955
rect 566 1912 572 1921
rect 624 1912 630 1964
rect 872 1964 924 1970
rect 715 1921 872 1955
rect 663 1906 715 1912
rect 1859 1968 1919 1977
rect 1829 1921 1859 1955
rect 872 1906 924 1912
rect 2759 1968 2819 1977
rect 2729 1921 2759 1955
rect 1859 1899 1919 1908
rect 2759 1899 2819 1908
rect 963 1603 1015 1609
rect 1259 1607 1319 1616
rect 1015 1560 1259 1594
rect 963 1545 1015 1551
rect 1259 1538 1319 1547
rect 509 1437 569 1446
rect 509 1368 569 1377
rect 1109 1437 1169 1446
rect 1109 1368 1169 1377
rect 1709 1437 1769 1446
rect 1709 1368 1769 1377
rect 2309 1437 2369 1446
rect 2309 1368 2369 1377
rect 209 1227 269 1236
rect 209 1158 269 1167
rect 809 1227 869 1236
rect 809 1158 869 1167
rect 1409 1227 1469 1236
rect 1409 1158 1469 1167
rect 2009 1227 2069 1236
rect 2009 1158 2069 1167
rect 2609 1227 2669 1236
rect 2609 1158 2669 1167
rect 359 1057 419 1066
rect 1772 1053 1824 1059
rect 419 1010 1772 1044
rect 359 988 419 997
rect 2672 1053 2724 1059
rect 1824 1010 2672 1044
rect 1772 995 1824 1001
rect 2672 995 2724 1001
rect 959 973 1019 982
rect 1472 969 1524 975
rect 1019 926 1472 960
rect 959 904 1019 913
rect 1472 911 1524 917
rect 659 889 719 898
rect 2372 885 2424 891
rect 719 842 2372 876
rect 659 820 719 829
rect 2372 827 2424 833
rect 1172 805 1224 807
rect 1172 801 1259 805
rect 972 758 1172 792
rect 1224 749 1259 801
rect 1172 745 1259 749
rect 1319 792 1328 805
rect 2072 801 2124 807
rect 1319 758 2072 792
rect 1319 745 1328 758
rect 1172 743 1224 745
rect 2072 743 2124 749
rect 663 622 715 628
rect 566 613 572 622
rect 148 579 572 613
rect 566 570 572 579
rect 624 570 630 622
rect 872 622 924 628
rect 715 579 872 613
rect 663 564 715 570
rect 1859 626 1919 635
rect 1829 579 1859 613
rect 872 564 924 570
rect 2759 626 2819 635
rect 2729 579 2759 613
rect 1859 557 1919 566
rect 2759 557 2819 566
rect 272 261 324 267
rect 148 218 272 252
rect 272 203 324 209
rect 509 95 569 104
rect 509 26 569 35
rect 1109 95 1169 104
rect 1109 26 1169 35
rect 1709 95 1769 104
rect 1709 26 1769 35
rect 2309 95 2369 104
rect 2309 26 2369 35
<< via2 >>
rect 209 2509 269 2569
rect 809 2509 869 2569
rect 1409 2509 1469 2569
rect 2009 2509 2069 2569
rect 2609 2509 2669 2569
rect 359 2339 419 2399
rect 959 2255 1019 2315
rect 659 2171 719 2231
rect 1859 1908 1919 1968
rect 2759 1908 2819 1968
rect 1259 1547 1319 1607
rect 509 1377 569 1437
rect 1109 1377 1169 1437
rect 1709 1377 1769 1437
rect 2309 1377 2369 1437
rect 209 1167 269 1227
rect 809 1167 869 1227
rect 1409 1167 1469 1227
rect 2009 1167 2069 1227
rect 2609 1167 2669 1227
rect 359 1053 419 1057
rect 359 1001 363 1053
rect 363 1001 415 1053
rect 415 1001 419 1053
rect 359 997 419 1001
rect 959 969 1019 973
rect 959 917 963 969
rect 963 917 1015 969
rect 1015 917 1019 969
rect 959 913 1019 917
rect 659 885 719 889
rect 659 833 663 885
rect 663 833 715 885
rect 715 833 719 885
rect 659 829 719 833
rect 1259 745 1319 805
rect 1859 566 1919 626
rect 2759 566 2819 626
rect 509 35 569 95
rect 1109 35 1169 95
rect 1709 35 1769 95
rect 2309 35 2369 95
<< metal3 >>
rect 204 2569 274 2574
rect 204 2509 209 2569
rect 269 2509 274 2569
rect 804 2569 874 2574
rect 204 2504 274 2509
rect 209 1232 269 2504
rect 354 2399 424 2404
rect 354 2339 359 2399
rect 419 2339 424 2399
rect 354 2334 424 2339
rect 204 1227 274 1232
rect 204 1167 209 1227
rect 269 1167 274 1227
rect 204 1162 274 1167
rect 209 36 269 1162
rect 359 1062 419 2334
rect 509 1442 569 2568
rect 804 2509 809 2569
rect 869 2509 874 2569
rect 1404 2569 1474 2574
rect 804 2504 874 2509
rect 654 2231 724 2236
rect 654 2171 659 2231
rect 719 2171 724 2231
rect 654 2166 724 2171
rect 504 1437 574 1442
rect 504 1377 509 1437
rect 569 1377 574 1437
rect 504 1372 574 1377
rect 354 1057 424 1062
rect 354 997 359 1057
rect 419 997 424 1057
rect 354 992 424 997
rect 509 100 569 1372
rect 659 894 719 2166
rect 809 1232 869 2504
rect 954 2315 1024 2320
rect 954 2255 959 2315
rect 1019 2255 1024 2315
rect 954 2250 1024 2255
rect 804 1227 874 1232
rect 804 1167 809 1227
rect 869 1167 874 1227
rect 804 1162 874 1167
rect 654 889 724 894
rect 654 829 659 889
rect 719 829 724 889
rect 654 824 724 829
rect 504 95 574 100
rect 504 35 509 95
rect 569 35 574 95
rect 809 36 869 1162
rect 959 978 1019 2250
rect 1109 1442 1169 2568
rect 1404 2509 1409 2569
rect 1469 2509 1474 2569
rect 2004 2569 2074 2574
rect 1404 2504 1474 2509
rect 1254 1607 1324 1612
rect 1254 1547 1259 1607
rect 1319 1547 1324 1607
rect 1254 1542 1324 1547
rect 1104 1437 1174 1442
rect 1104 1377 1109 1437
rect 1169 1377 1174 1437
rect 1104 1372 1174 1377
rect 954 973 1024 978
rect 954 913 959 973
rect 1019 913 1024 973
rect 954 908 1024 913
rect 1109 100 1169 1372
rect 1259 810 1319 1542
rect 1409 1232 1469 2504
rect 1709 1442 1769 2568
rect 2004 2509 2009 2569
rect 2069 2509 2074 2569
rect 2604 2569 2674 2574
rect 2004 2504 2074 2509
rect 1859 1973 1919 2072
rect 1854 1968 1924 1973
rect 1854 1908 1859 1968
rect 1919 1908 1924 1968
rect 1854 1903 1924 1908
rect 1859 1804 1919 1903
rect 1704 1437 1774 1442
rect 1704 1377 1709 1437
rect 1769 1377 1774 1437
rect 1704 1372 1774 1377
rect 1404 1227 1474 1232
rect 1404 1167 1409 1227
rect 1469 1167 1474 1227
rect 1404 1162 1474 1167
rect 1254 805 1324 810
rect 1254 745 1259 805
rect 1319 745 1324 805
rect 1254 740 1324 745
rect 1104 95 1174 100
rect 504 30 574 35
rect 1104 35 1109 95
rect 1169 35 1174 95
rect 1409 36 1469 1162
rect 1709 100 1769 1372
rect 2009 1232 2069 2504
rect 2309 1442 2369 2568
rect 2604 2509 2609 2569
rect 2669 2509 2674 2569
rect 2604 2504 2674 2509
rect 2304 1437 2374 1442
rect 2304 1377 2309 1437
rect 2369 1377 2374 1437
rect 2304 1372 2374 1377
rect 2004 1227 2074 1232
rect 2004 1167 2009 1227
rect 2069 1167 2074 1227
rect 2004 1162 2074 1167
rect 1859 631 1919 730
rect 1854 626 1924 631
rect 1854 566 1859 626
rect 1919 566 1924 626
rect 1854 561 1924 566
rect 1859 462 1919 561
rect 1704 95 1774 100
rect 1104 30 1174 35
rect 1704 35 1709 95
rect 1769 35 1774 95
rect 2009 36 2069 1162
rect 2309 100 2369 1372
rect 2609 1232 2669 2504
rect 2759 1973 2819 2072
rect 2754 1968 2824 1973
rect 2754 1908 2759 1968
rect 2819 1908 2824 1968
rect 2754 1903 2824 1908
rect 2759 1804 2819 1903
rect 2604 1227 2674 1232
rect 2604 1167 2609 1227
rect 2669 1167 2674 1227
rect 2604 1162 2674 1167
rect 2304 95 2374 100
rect 1704 30 1774 35
rect 2304 35 2309 95
rect 2369 35 2374 95
rect 2609 36 2669 1162
rect 2759 631 2819 730
rect 2754 626 2824 631
rect 2754 566 2759 626
rect 2819 566 2824 626
rect 2754 561 2824 566
rect 2759 462 2819 561
rect 2304 30 2374 35
use transistor_pair_bus9  transistor_pair_bus9_0
timestamp 1727641816
transform 1 0 60 0 1 0
box -60 0 2936 1292
use transistor_pair_bus9  transistor_pair_bus9_1
timestamp 1727641816
transform 1 0 60 0 1 1342
box -60 0 2936 1292
use inverter  x1
timestamp 1727638268
transform 1 0 60 0 1 0
box 88 36 388 1226
use inverter  x2
timestamp 1727638268
transform 1 0 360 0 1 0
box 88 36 388 1226
use inverter  x3
timestamp 1727638268
transform 1 0 660 0 1 0
box 88 36 388 1226
use inverter  x4
timestamp 1727638268
transform 1 0 360 0 1 1342
box 88 36 388 1226
use inverter  x5
timestamp 1727638268
transform 1 0 660 0 1 1342
box 88 36 388 1226
use nor3  x6
timestamp 1727641975
transform 1 0 960 0 1 0
box 88 36 964 1226
use nor3  x7
timestamp 1727641975
transform 1 0 1860 0 1 0
box 88 36 964 1226
use nor3  x8
timestamp 1727641975
transform 1 0 960 0 1 1342
box 88 36 964 1226
use nor3  x9
timestamp 1727641975
transform 1 0 1860 0 1 1342
box 88 36 964 1226
use inverter  xdummy
timestamp 1727638268
transform 1 0 60 0 1 1342
box 88 36 388 1226
<< labels >>
flabel metal2 148 218 272 252 0 FreeSans 128 0 0 0 EN
port 2 nsew
flabel metal2 148 579 572 613 0 FreeSans 128 0 0 0 D0
port 0 nsew
flabel metal2 148 1921 572 1955 0 FreeSans 128 0 0 0 D1
port 1 nsew
flabel metal3 1859 462 1919 730 0 FreeSans 128 0 0 0 U0
port 3 nsew
flabel metal3 2759 462 2819 730 0 FreeSans 128 0 0 0 U1
port 4 nsew
flabel metal3 1859 1804 1919 2072 0 FreeSans 128 0 0 0 U2
port 5 nsew
flabel metal3 2759 1804 2819 2072 0 FreeSans 128 0 0 0 U3
port 6 nsew
flabel metal3 209 36 269 2568 0 FreeSans 128 0 0 0 VDD
port 7 nsew
flabel metal3 509 36 569 2568 0 FreeSans 128 0 0 0 VSS
port 8 nsew
<< end >>
