magic
tech sky130A
magscale 1 2
timestamp 1727641773
<< metal1 >>
rect 2268 9347 2328 9353
rect 2600 9347 2660 9353
rect 2932 9347 2992 9353
rect 3264 9347 3324 9353
rect 3596 9347 3656 9353
rect 3928 9347 3988 9353
rect 276 8915 512 9347
rect 608 8915 844 9347
rect 940 8915 1176 9347
rect 1272 8915 1508 9347
rect 1604 9139 1840 9347
rect 1664 9079 1840 9139
rect 1604 8915 1840 9079
rect 1936 9264 2172 9347
rect 1996 9204 2172 9264
rect 1936 8915 2172 9204
rect 2328 9287 2504 9347
rect 2268 8915 2504 9287
rect 2660 9287 2836 9347
rect 2600 8915 2836 9287
rect 2992 9287 3168 9347
rect 2932 8915 3168 9287
rect 3324 9287 3500 9347
rect 3264 8915 3500 9287
rect 3656 9287 3832 9347
rect 3596 8915 3832 9287
rect 3988 9287 4164 9347
rect 3928 8915 4164 9287
rect 1438 2825 1498 2831
rect 1438 2547 1498 2765
rect 1770 2700 1830 2706
rect 1770 2547 1830 2640
rect 2102 2575 2162 2581
rect 276 2115 346 2547
rect 442 2115 678 2547
rect 774 2115 1010 2547
rect 1106 2115 1342 2547
rect 1438 2115 1674 2547
rect 1770 2115 2006 2547
rect 2162 2515 2338 2547
rect 2102 2115 2338 2515
rect 2434 2450 2670 2547
rect 2494 2390 2670 2450
rect 2434 2115 2670 2390
rect 2766 2325 3002 2547
rect 2826 2265 3002 2325
rect 2766 2115 3002 2265
rect 3098 2200 3334 2547
rect 3158 2140 3334 2200
rect 3098 2115 3334 2140
rect 3430 2115 3666 2547
rect 3762 2115 3998 2547
rect 3430 2075 3490 2115
rect 3430 2009 3490 2015
rect 3304 1950 3364 1956
rect 3762 1950 3822 2115
rect 3298 1890 3304 1950
rect 3364 1890 3822 1950
rect 3304 1884 3364 1890
rect 3430 1825 3490 1831
rect 4099 1825 4159 2547
rect 3424 1765 3430 1825
rect 3490 1765 4159 1825
rect 3430 1759 3490 1765
<< via1 >>
rect 1604 9079 1664 9139
rect 1936 9204 1996 9264
rect 2268 9287 2328 9347
rect 2600 9287 2660 9347
rect 2932 9287 2992 9347
rect 3264 9287 3324 9347
rect 3596 9287 3656 9347
rect 3928 9287 3988 9347
rect 1438 2765 1498 2825
rect 1770 2640 1830 2700
rect 2102 2515 2162 2575
rect 2434 2390 2494 2450
rect 2766 2265 2826 2325
rect 3098 2140 3158 2200
rect 3430 2015 3490 2075
rect 3304 1890 3364 1950
rect 3430 1765 3490 1825
<< metal2 >>
rect 277 11273 415 11411
rect 665 10988 783 10998
rect 665 10890 675 10988
rect 773 10890 783 10988
rect 665 10880 783 10890
rect 941 10988 1059 10998
rect 941 10890 951 10988
rect 1049 10890 1059 10988
rect 941 10880 1059 10890
rect 1217 10988 1335 10998
rect 1217 10890 1227 10988
rect 1325 10890 1335 10988
rect 1217 10880 1335 10890
rect 1493 10988 1611 10998
rect 1493 10890 1503 10988
rect 1601 10890 1611 10988
rect 1493 10880 1611 10890
rect 1769 10988 1887 10998
rect 1769 10890 1779 10988
rect 1877 10890 1887 10988
rect 1769 10880 1887 10890
rect 2045 10988 2163 10998
rect 2045 10890 2055 10988
rect 2153 10890 2163 10988
rect 2045 10880 2163 10890
rect 2321 10988 2439 10998
rect 2321 10890 2331 10988
rect 2429 10890 2439 10988
rect 2321 10880 2439 10890
rect 2597 10988 2715 10998
rect 2597 10890 2607 10988
rect 2705 10890 2715 10988
rect 2597 10880 2715 10890
rect 2268 9347 2328 9356
rect 2600 9347 2660 9356
rect 2932 9347 2992 9356
rect 3264 9347 3324 9356
rect 3596 9347 3656 9356
rect 3928 9347 3988 9356
rect 2262 9287 2268 9347
rect 2328 9287 2334 9347
rect 2594 9287 2600 9347
rect 2660 9287 2666 9347
rect 2926 9287 2932 9347
rect 2992 9287 2998 9347
rect 3258 9287 3264 9347
rect 3324 9287 3330 9347
rect 3590 9287 3596 9347
rect 3656 9287 3662 9347
rect 3922 9287 3928 9347
rect 3988 9287 3994 9347
rect 2268 9278 2328 9287
rect 2600 9278 2660 9287
rect 2932 9278 2992 9287
rect 3264 9278 3324 9287
rect 3596 9278 3656 9287
rect 3928 9278 3988 9287
rect 1936 9264 1996 9273
rect 1930 9204 1936 9264
rect 1996 9204 2002 9264
rect 1936 9195 1996 9204
rect 1604 9139 1664 9148
rect 1598 9079 1604 9139
rect 1664 9079 1670 9139
rect 1604 9070 1664 9079
rect 1438 2825 1498 2834
rect 1432 2765 1438 2825
rect 1498 2765 1504 2825
rect 1438 2756 1498 2765
rect 1770 2700 1830 2709
rect 1764 2640 1770 2700
rect 1830 2640 1836 2700
rect 1770 2631 1830 2640
rect 2102 2575 2162 2584
rect 2096 2515 2102 2575
rect 2162 2515 2168 2575
rect 2102 2506 2162 2515
rect 2434 2450 2494 2459
rect 2434 2381 2494 2390
rect 2766 2325 2826 2334
rect 2760 2265 2766 2325
rect 2826 2265 2832 2325
rect 2766 2256 2826 2265
rect 3098 2200 3158 2209
rect 3092 2140 3098 2200
rect 3158 2140 3164 2200
rect 3098 2131 3158 2140
rect 3430 2075 3490 2084
rect 3424 2015 3430 2075
rect 3490 2015 3496 2075
rect 3430 2006 3490 2015
rect 3304 1950 3364 1959
rect 3298 1890 3304 1950
rect 3364 1890 3370 1950
rect 3304 1881 3364 1890
rect 3430 1825 3490 1831
rect 3421 1765 3430 1825
rect 3490 1765 3499 1825
rect 3430 1759 3490 1765
rect 562 557 680 675
rect 552 493 690 513
rect 552 395 572 493
rect 670 395 690 493
rect 552 375 690 395
rect 838 493 956 503
rect 838 395 848 493
rect 946 395 956 493
rect 838 385 956 395
rect 1114 493 1232 503
rect 1114 395 1124 493
rect 1222 395 1232 493
rect 1114 385 1232 395
rect 1390 493 1508 503
rect 1390 395 1400 493
rect 1498 395 1508 493
rect 1390 385 1508 395
rect 1666 493 1784 503
rect 1666 395 1676 493
rect 1774 395 1784 493
rect 1666 385 1784 395
rect 1942 493 2060 503
rect 1942 395 1952 493
rect 2050 395 2060 493
rect 1942 385 2060 395
rect 2218 493 2336 503
rect 2218 395 2228 493
rect 2326 395 2336 493
rect 2218 385 2336 395
rect 2494 493 2612 503
rect 2494 395 2504 493
rect 2602 395 2612 493
rect 2494 385 2612 395
rect 276 42 414 180
<< via2 >>
rect 675 10890 773 10988
rect 951 10890 1049 10988
rect 1227 10890 1325 10988
rect 1503 10890 1601 10988
rect 1779 10890 1877 10988
rect 2055 10890 2153 10988
rect 2331 10890 2429 10988
rect 2607 10890 2705 10988
rect 563 9964 681 10082
rect 839 9964 957 10082
rect 1115 9964 1233 10082
rect 1391 9964 1509 10082
rect 1667 9964 1785 10082
rect 1943 9964 2061 10082
rect 2219 9964 2337 10082
rect 2495 9964 2613 10082
rect 2268 9287 2328 9347
rect 2600 9287 2660 9347
rect 2932 9287 2992 9347
rect 3264 9287 3324 9347
rect 3596 9287 3656 9347
rect 3928 9287 3988 9347
rect 1936 9204 1996 9264
rect 1604 9079 1664 9139
rect 1438 2765 1498 2825
rect 1770 2640 1830 2700
rect 2102 2515 2162 2575
rect 2434 2390 2494 2450
rect 2766 2265 2826 2325
rect 3098 2140 3158 2200
rect 3430 2015 3490 2075
rect 3304 1890 3364 1950
rect 562 1660 680 1778
rect 838 1659 956 1777
rect 1114 1659 1232 1777
rect 1390 1659 1508 1777
rect 1666 1659 1784 1777
rect 1942 1659 2060 1777
rect 2218 1659 2336 1777
rect 2494 1659 2612 1777
rect 3430 1765 3490 1825
rect 572 395 670 493
rect 848 395 946 493
rect 1124 395 1222 493
rect 1400 395 1498 493
rect 1676 395 1774 493
rect 1952 395 2050 493
rect 2228 395 2326 493
rect 2504 395 2602 493
<< metal3 >>
rect 665 10988 783 10998
rect 665 10890 675 10988
rect 773 10890 783 10988
rect 665 10880 783 10890
rect 941 10988 1059 10998
rect 941 10890 951 10988
rect 1049 10890 1059 10988
rect 941 10880 1059 10890
rect 1217 10988 1335 10998
rect 1217 10890 1227 10988
rect 1325 10890 1335 10988
rect 1217 10880 1335 10890
rect 1493 10988 1611 10998
rect 1493 10890 1503 10988
rect 1601 10890 1611 10988
rect 1493 10880 1611 10890
rect 1769 10988 1887 10998
rect 1769 10890 1779 10988
rect 1877 10890 1887 10988
rect 1769 10880 1887 10890
rect 2045 10988 2163 10998
rect 2045 10890 2055 10988
rect 2153 10890 2163 10988
rect 2045 10880 2163 10890
rect 2321 10988 2439 10998
rect 2321 10890 2331 10988
rect 2429 10890 2439 10988
rect 2321 10880 2439 10890
rect 2597 10988 2715 10998
rect 2597 10890 2607 10988
rect 2705 10890 2715 10988
rect 2597 10880 2715 10890
rect 138 10600 793 10738
rect 138 1331 276 10600
rect 553 10082 691 10092
rect 553 9964 563 10082
rect 681 9964 691 10082
rect 553 9954 691 9964
rect 829 10082 967 10092
rect 829 9964 839 10082
rect 957 9964 967 10082
rect 829 9954 967 9964
rect 1105 10082 1243 10092
rect 1105 9964 1115 10082
rect 1233 9964 1243 10082
rect 1105 9954 1243 9964
rect 1381 10082 1519 10092
rect 1381 9964 1391 10082
rect 1509 9964 1519 10082
rect 1381 9954 1519 9964
rect 1657 10082 1795 10092
rect 1657 9964 1667 10082
rect 1785 9964 1795 10082
rect 1657 9954 1795 9964
rect 1933 10082 2071 10092
rect 1933 9964 1943 10082
rect 2061 9964 2071 10082
rect 1933 9954 2071 9964
rect 2209 10082 2347 10092
rect 2209 9964 2219 10082
rect 2337 9964 2347 10082
rect 2209 9954 2347 9964
rect 2485 10082 2623 10092
rect 2485 9964 2495 10082
rect 2613 10014 2623 10082
rect 2613 9964 3988 10014
rect 2485 9954 3988 9964
rect 631 9139 691 9954
rect 907 9264 967 9954
rect 1183 9389 1243 9954
rect 1459 9514 1519 9954
rect 1735 9639 1795 9954
rect 2011 9764 2071 9954
rect 2287 9889 2347 9954
rect 2287 9829 3656 9889
rect 2011 9704 3324 9764
rect 1735 9579 2992 9639
rect 1459 9454 2660 9514
rect 1183 9352 2328 9389
rect 2600 9352 2660 9454
rect 2932 9352 2992 9579
rect 3264 9352 3324 9704
rect 3596 9352 3656 9829
rect 3928 9352 3988 9954
rect 1183 9347 2333 9352
rect 1183 9329 2268 9347
rect 2263 9287 2268 9329
rect 2328 9287 2333 9347
rect 2263 9282 2333 9287
rect 2595 9347 2665 9352
rect 2595 9287 2600 9347
rect 2660 9287 2665 9347
rect 2595 9282 2665 9287
rect 2927 9347 2997 9352
rect 2927 9287 2932 9347
rect 2992 9287 2997 9347
rect 2927 9282 2997 9287
rect 3259 9347 3329 9352
rect 3259 9287 3264 9347
rect 3324 9287 3329 9347
rect 3259 9282 3329 9287
rect 3591 9347 3661 9352
rect 3591 9287 3596 9347
rect 3656 9287 3661 9347
rect 3591 9282 3661 9287
rect 3923 9347 3993 9352
rect 3923 9287 3928 9347
rect 3988 9287 3993 9347
rect 3923 9282 3993 9287
rect 1931 9264 2001 9269
rect 907 9204 1936 9264
rect 1996 9204 2001 9264
rect 1931 9199 2001 9204
rect 1599 9139 1669 9144
rect 631 9079 1604 9139
rect 1664 9079 1669 9139
rect 1599 9074 1669 9079
rect 1433 2825 1503 2830
rect 630 2765 1438 2825
rect 1498 2765 1503 2825
rect 630 1788 690 2765
rect 1433 2760 1503 2765
rect 1765 2700 1835 2705
rect 552 1778 690 1788
rect 906 2640 1770 2700
rect 1830 2640 1835 2700
rect 906 1787 966 2640
rect 1765 2635 1835 2640
rect 2097 2575 2167 2580
rect 1182 2515 2102 2575
rect 2162 2515 2167 2575
rect 1182 1787 1242 2515
rect 2097 2510 2167 2515
rect 2429 2450 2499 2455
rect 1458 2390 2434 2450
rect 2494 2390 2499 2450
rect 1458 1787 1518 2390
rect 2429 2385 2499 2390
rect 2761 2325 2831 2330
rect 1734 2265 2766 2325
rect 2826 2265 2831 2325
rect 1734 1787 1794 2265
rect 2761 2260 2831 2265
rect 3093 2200 3163 2205
rect 2010 2140 3098 2200
rect 3158 2140 3163 2200
rect 2010 1787 2070 2140
rect 3093 2135 3163 2140
rect 3425 2075 3495 2080
rect 2286 2015 3430 2075
rect 3490 2015 3495 2075
rect 2286 1787 2346 2015
rect 3425 2010 3495 2015
rect 3299 1950 3369 1955
rect 2562 1890 3304 1950
rect 3364 1890 3369 1950
rect 2562 1787 2622 1890
rect 3299 1885 3369 1890
rect 3425 1825 3495 1830
rect 2838 1787 3430 1825
rect 552 1660 562 1778
rect 680 1660 690 1778
rect 552 1650 690 1660
rect 828 1777 966 1787
rect 828 1659 838 1777
rect 956 1659 966 1777
rect 828 1649 966 1659
rect 1104 1777 1242 1787
rect 1104 1659 1114 1777
rect 1232 1659 1242 1777
rect 1104 1649 1242 1659
rect 1380 1777 1518 1787
rect 1380 1659 1390 1777
rect 1508 1659 1518 1777
rect 1380 1649 1518 1659
rect 1656 1777 1794 1787
rect 1656 1659 1666 1777
rect 1784 1659 1794 1777
rect 1656 1649 1794 1659
rect 1932 1777 2070 1787
rect 1932 1659 1942 1777
rect 2060 1659 2070 1777
rect 1932 1649 2070 1659
rect 2208 1777 2346 1787
rect 2208 1659 2218 1777
rect 2336 1659 2346 1777
rect 2208 1649 2346 1659
rect 2484 1777 2622 1787
rect 2484 1659 2494 1777
rect 2612 1659 2622 1777
rect 2484 1649 2622 1659
rect 2760 1765 3430 1787
rect 3490 1765 3495 1825
rect 2760 1649 2898 1765
rect 3425 1760 3495 1765
rect 138 1193 792 1331
rect 562 493 680 503
rect 562 395 572 493
rect 670 395 680 493
rect 562 385 680 395
rect 838 493 956 503
rect 838 395 848 493
rect 946 395 956 493
rect 838 385 956 395
rect 1114 493 1232 503
rect 1114 395 1124 493
rect 1222 395 1232 493
rect 1114 385 1232 395
rect 1390 493 1508 503
rect 1390 395 1400 493
rect 1498 395 1508 493
rect 1390 385 1508 395
rect 1666 493 1784 503
rect 1666 395 1676 493
rect 1774 395 1784 493
rect 1666 385 1784 395
rect 1942 493 2060 503
rect 1942 395 1952 493
rect 2050 395 2060 493
rect 1942 385 2060 395
rect 2218 493 2336 503
rect 2218 395 2228 493
rect 2326 395 2336 493
rect 2218 385 2336 395
rect 2494 493 2612 503
rect 2494 395 2504 493
rect 2602 395 2612 493
rect 2494 385 2612 395
use passgates  passgates_0
timestamp 1727641178
transform 1 0 111 0 1 9407
box 0 0 3056 2076
use passgates  passgates_1
timestamp 1727641178
transform 1 0 110 0 1 0
box 0 0 3056 2076
use sky130_fd_pr__res_xhigh_po_0p35_EMC64D  sky130_fd_pr__res_xhigh_po_0p35_EMC64D_0
timestamp 1727597281
transform 1 0 2220 0 1 5731
box -2110 -3616 2110 3616
<< labels >>
flabel metal3 665 10880 783 10998 0 FreeSans 128 0 0 0 U1
port 3 nsew
flabel metal3 941 10880 1059 10998 0 FreeSans 128 0 0 0 U3
port 5 nsew
flabel metal3 1217 10880 1335 10998 0 FreeSans 128 0 0 0 U5
port 7 nsew
flabel metal3 1493 10880 1611 10998 0 FreeSans 128 0 0 0 U7
port 9 nsew
flabel metal3 1769 10880 1887 10998 0 FreeSans 128 0 0 0 U9
port 11 nsew
flabel metal3 2045 10880 2163 10998 0 FreeSans 128 0 0 0 U11
port 13 nsew
flabel metal3 2321 10880 2439 10998 0 FreeSans 128 0 0 0 U13
port 15 nsew
flabel metal3 2597 10880 2715 10998 0 FreeSans 128 0 0 0 U15
port 17 nsew
flabel metal3 2760 1649 2898 1787 0 FreeSans 128 0 0 0 B
port 1 nsew
flabel metal3 552 1650 690 1788 0 FreeSans 128 0 0 0 A
port 0 nsew
flabel metal3 654 1193 792 1331 0 FreeSans 128 0 0 0 W
port 20 nsew
flabel metal2 276 42 414 180 0 FreeSans 128 0 0 0 VSS
port 19 nsew
flabel metal3 562 385 680 503 0 FreeSans 128 0 0 0 U0
port 2 nsew
flabel metal3 2494 385 2612 503 0 FreeSans 128 0 0 0 U14
port 16 nsew
flabel metal3 2218 385 2336 503 0 FreeSans 128 0 0 0 U12
port 14 nsew
flabel metal3 1942 385 2060 503 0 FreeSans 128 0 0 0 U10
port 12 nsew
flabel metal3 1666 385 1784 503 0 FreeSans 128 0 0 0 U8
port 10 nsew
flabel metal3 1390 385 1508 503 0 FreeSans 128 0 0 0 U6
port 8 nsew
flabel metal3 1114 385 1232 503 0 FreeSans 128 0 0 0 U4
port 6 nsew
flabel metal3 838 385 956 503 0 FreeSans 128 0 0 0 U2
port 4 nsew
flabel metal2 277 11273 415 11411 0 FreeSans 128 0 0 0 VDD
port 18 nsew
<< end >>
