magic
tech sky130A
magscale 1 2
timestamp 1727607772
<< metal1 >>
rect 3074 11099 3212 11105
rect 3212 10961 7274 11099
rect 3074 10955 3212 10961
rect 3074 9887 3212 9893
rect 3212 9749 7274 9887
rect 3074 9743 3212 9749
rect 3074 1705 3212 1711
rect 3212 1567 7274 1705
rect 3074 1561 3212 1567
rect 3074 493 3212 499
rect 3212 355 7274 493
rect 3074 349 3212 355
<< via1 >>
rect 3074 10961 3212 11099
rect 3074 9749 3212 9887
rect 3074 1567 3212 1705
rect 3074 355 3212 493
<< metal2 >>
rect 4504 11874 4538 12445
rect 4364 11840 4538 11874
rect 4225 11622 4285 11631
rect 4364 11609 4398 11840
rect 4285 11575 4398 11609
rect 4490 11714 4550 11748
rect 4225 11553 4285 11562
rect 4099 11496 4159 11505
rect 4490 11483 4524 11714
rect 4159 11449 4524 11483
rect 4099 11427 4159 11436
rect 277 11273 415 11411
rect 2761 11273 3212 11411
rect 3074 11099 3212 11273
rect 4477 11116 4537 11125
rect 3068 10961 3074 11099
rect 3212 10961 3218 11099
rect 4477 11047 4537 11056
rect 4351 10419 4411 10428
rect 4411 10372 4538 10406
rect 4351 10350 4411 10359
rect 3973 10293 4033 10302
rect 4477 10293 4537 10302
rect 4033 10246 4477 10280
rect 3973 10224 4033 10233
rect 4477 10224 4537 10233
rect 3847 10167 3907 10176
rect 4351 10167 4411 10176
rect 3907 10120 4351 10154
rect 3847 10098 3907 10107
rect 4351 10098 4411 10107
rect 3068 9749 3074 9887
rect 3212 9749 3218 9887
rect 4477 9774 4537 9783
rect 3074 9587 3212 9749
rect 4477 9705 4537 9714
rect 2761 9449 3212 9587
rect 4351 9077 4411 9086
rect 4411 9030 4538 9064
rect 4351 9008 4411 9017
rect 4225 8432 4285 8441
rect 4285 8385 4538 8419
rect 4225 8363 4285 8372
rect 4099 7735 4159 7744
rect 4159 7688 4538 7722
rect 4099 7666 4159 7675
rect 3595 7090 3655 7099
rect 3655 7043 4538 7077
rect 3595 7021 3655 7030
rect 3721 6393 3781 6402
rect 3781 6346 4538 6380
rect 3721 6324 3781 6333
rect 4477 5748 4537 5757
rect 4477 5679 4537 5688
rect 4351 5051 4411 5060
rect 4411 5004 4538 5038
rect 4351 4982 4411 4991
rect 4099 4406 4159 4415
rect 4159 4359 4538 4393
rect 4099 4337 4159 4346
rect 4225 3709 4285 3718
rect 4285 3662 4538 3696
rect 6850 3662 7727 3696
rect 4225 3640 4285 3649
rect 3847 3064 3907 3073
rect 3907 3017 4538 3051
rect 3847 2995 3907 3004
rect 3973 2367 4033 2376
rect 4033 2320 4538 2354
rect 6850 2320 7727 2354
rect 3973 2298 4033 2307
rect 2760 1866 3212 2004
rect 3074 1705 3212 1866
rect 3068 1567 3074 1705
rect 3212 1567 3218 1705
rect 6850 978 7727 1012
rect 3068 355 3074 493
rect 3212 355 3218 493
rect 3074 180 3212 355
rect 276 42 414 180
rect 2760 42 3212 180
rect 6850 -364 7727 -330
<< via2 >>
rect 4225 11562 4285 11622
rect 4099 11436 4159 11496
rect 4477 11056 4537 11116
rect 4351 10359 4411 10419
rect 3973 10233 4033 10293
rect 4477 10233 4537 10293
rect 3847 10107 3907 10167
rect 4351 10107 4411 10167
rect 4477 9714 4537 9774
rect 4351 9017 4411 9077
rect 4225 8372 4285 8432
rect 4099 7675 4159 7735
rect 3595 7030 3655 7090
rect 3721 6333 3781 6393
rect 4477 5688 4537 5748
rect 4351 4991 4411 5051
rect 4099 4346 4159 4406
rect 4225 3649 4285 3709
rect 3847 3004 3907 3064
rect 3973 2307 4033 2367
rect 562 569 680 679
<< metal3 >>
rect 694 11814 4537 11874
rect 694 10909 754 11814
rect 970 11688 4411 11748
rect 970 10909 1030 11688
rect 4220 11622 4290 11627
rect 1246 11562 4225 11622
rect 4285 11562 4290 11622
rect 1246 10909 1306 11562
rect 4220 11557 4290 11562
rect 4094 11496 4164 11501
rect 1522 11436 4099 11496
rect 4159 11436 4164 11496
rect 1522 10909 1582 11436
rect 4094 11431 4164 11436
rect 1798 11310 4285 11370
rect 1798 10909 1858 11310
rect 2074 11184 4159 11244
rect 2074 10909 2134 11184
rect 2350 11058 4033 11118
rect 2350 10909 2410 11058
rect 2626 10909 3907 10969
rect 3847 10172 3907 10909
rect 3973 10298 4033 11058
rect 3968 10293 4038 10298
rect 3968 10233 3973 10293
rect 4033 10233 4038 10293
rect 3968 10228 4038 10233
rect 3842 10167 3912 10172
rect 3842 10107 3847 10167
rect 3907 10107 3912 10167
rect 3842 10102 3912 10107
rect 4099 7740 4159 11184
rect 4225 8437 4285 11310
rect 4351 10424 4411 11688
rect 4477 11121 4537 11814
rect 4472 11116 4542 11121
rect 4472 11056 4477 11116
rect 4537 11056 4542 11116
rect 4472 11051 4542 11056
rect 4346 10419 4416 10424
rect 4346 10359 4351 10419
rect 4411 10359 4416 10419
rect 4346 10354 4416 10359
rect 4472 10293 4542 10298
rect 4472 10233 4477 10293
rect 4537 10233 4542 10293
rect 4472 10228 4542 10233
rect 4346 10167 4416 10172
rect 4346 10107 4351 10167
rect 4411 10107 4416 10167
rect 4346 10102 4416 10107
rect 4351 9082 4411 10102
rect 4477 9779 4537 10228
rect 4472 9774 4542 9779
rect 4472 9714 4477 9774
rect 4537 9714 4542 9774
rect 4472 9709 4542 9714
rect 4346 9077 4416 9082
rect 4346 9017 4351 9077
rect 4411 9017 4416 9077
rect 4346 9012 4416 9017
rect 4220 8432 4290 8437
rect 4220 8372 4225 8432
rect 4285 8372 4290 8432
rect 4220 8367 4290 8372
rect 4094 7735 4164 7740
rect 4094 7675 4099 7735
rect 4159 7675 4164 7735
rect 4094 7670 4164 7675
rect 3590 7090 3660 7095
rect 3590 7030 3595 7090
rect 3655 7030 3660 7090
rect 3590 7025 3660 7030
rect 2760 1649 2898 1787
rect 654 1193 792 1331
rect 3595 1127 3655 7025
rect 3716 6393 3786 6398
rect 3716 6333 3721 6393
rect 3781 6333 3786 6393
rect 3716 6328 3786 6333
rect 1143 1067 3655 1127
rect 552 679 690 701
rect 552 569 562 679
rect 680 569 690 679
rect 552 563 690 569
rect 591 199 651 474
rect 867 325 927 474
rect 1143 414 1203 1067
rect 3721 1001 3781 6328
rect 4472 5748 4542 5753
rect 4472 5688 4477 5748
rect 4537 5688 4542 5748
rect 4472 5683 4542 5688
rect 4346 5051 4416 5056
rect 4346 4991 4351 5051
rect 4411 4991 4416 5051
rect 4346 4986 4416 4991
rect 4094 4406 4164 4411
rect 4094 4346 4099 4406
rect 4159 4346 4164 4406
rect 4094 4341 4164 4346
rect 3842 3064 3912 3069
rect 3842 3004 3847 3064
rect 3907 3004 3912 3064
rect 3842 2999 3912 3004
rect 1419 941 3781 1001
rect 1419 414 1479 941
rect 3847 875 3907 2999
rect 3968 2367 4038 2372
rect 3968 2307 3973 2367
rect 4033 2307 4038 2367
rect 3968 2302 4038 2307
rect 1695 815 3907 875
rect 1695 414 1755 815
rect 3973 749 4033 2302
rect 1971 689 4033 749
rect 1971 414 2031 689
rect 4099 623 4159 4341
rect 4220 3709 4290 3714
rect 4220 3649 4225 3709
rect 4285 3649 4290 3709
rect 4220 3644 4290 3649
rect 2247 563 4159 623
rect 2247 414 2307 563
rect 4225 474 4285 3644
rect 2523 414 4285 474
rect 4351 325 4411 4986
rect 867 265 4411 325
rect 4477 199 4537 5683
rect 591 139 4537 199
use decoder4_signed  decoder4_signed_0
timestamp 1727607772
transform -1 0 7422 0 1 -943
box -305 0 2996 13410
use digipot_1hot  x2
timestamp 1727597281
transform 1 0 0 0 1 0
box 110 0 4330 11483
<< labels >>
flabel metal2 276 42 414 180 0 FreeSans 128 0 0 0 VSS
port 7 nsew
flabel metal3 552 563 690 701 0 FreeSans 128 0 0 0 A
port 0 nsew
flabel metal3 2760 1649 2898 1787 0 FreeSans 128 0 0 0 B
port 1 nsew
flabel metal3 654 1193 792 1331 0 FreeSans 128 0 0 0 W
port 8 nsew
flabel metal2 6850 -364 7727 -330 0 FreeSans 128 0 0 0 D3
port 5 nsew
flabel metal2 6850 978 7727 1012 0 FreeSans 128 0 0 0 D0
port 2 nsew
flabel metal2 6850 2320 7727 2354 0 FreeSans 128 0 0 0 D1
port 3 nsew
flabel metal2 6850 3662 7727 3696 0 FreeSans 128 0 0 0 D2
port 4 nsew
flabel metal2 277 11273 415 11411 0 FreeSans 128 0 0 0 VDD
port 6 nsew
<< end >>
