magic
tech sky130A
magscale 1 2
timestamp 1727638502
use shifter_split  shifter_split_1
array 0 7 300 0 0 6127
timestamp 1727638502
transform 1 0 0 0 1 0
box 88 36 388 6061
use transistor_pair_bus8  transistor_pair_bus8_0
timestamp 1727637843
transform 1 0 0 0 1 0
box -60 0 2636 1292
use transistor_pair_bus8  transistor_pair_bus8_1
timestamp 1727637843
transform 1 0 0 0 1 1342
box -60 0 2636 1292
use transistor_pair_bus8  transistor_pair_bus8_2
timestamp 1727637843
transform 1 0 0 0 1 4835
box -60 0 2636 1292
<< end >>
