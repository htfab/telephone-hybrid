magic
tech sky130A
timestamp 1727635162
<< metal2 >>
rect 1400 2296 1792 2324
rect 1148 2268 2016 2296
rect 952 2240 2128 2268
rect 840 2212 2240 2240
rect 756 2184 2324 2212
rect 700 2156 2380 2184
rect 644 2128 2464 2156
rect 588 2100 2520 2128
rect 560 2072 2548 2100
rect 504 2044 2604 2072
rect 476 2016 2660 2044
rect 448 1988 2688 2016
rect 420 1960 1316 1988
rect 1848 1960 2716 1988
rect 420 1932 1148 1960
rect 2044 1932 2744 1960
rect 392 1904 1008 1932
rect 2128 1904 2772 1932
rect 364 1876 952 1904
rect 2212 1876 2772 1904
rect 364 1848 896 1876
rect 2240 1848 2800 1876
rect 364 1820 868 1848
rect 2268 1820 2800 1848
rect 336 1792 868 1820
rect 2296 1792 2800 1820
rect 336 1568 840 1792
rect 1064 1764 1232 1792
rect 1904 1764 2072 1792
rect 1008 1736 1260 1764
rect 1876 1736 2128 1764
rect 1008 1708 1288 1736
rect 1876 1708 2156 1736
rect 980 1680 1288 1708
rect 980 1624 1316 1680
rect 1848 1652 2156 1708
rect 1400 1624 1736 1652
rect 1820 1624 2156 1652
rect 1008 1568 2128 1624
rect 364 1540 840 1568
rect 364 1484 812 1540
rect 1036 1512 2128 1568
rect 2296 1568 2828 1792
rect 2296 1540 2800 1568
rect 2324 1512 2800 1540
rect 392 1456 756 1484
rect 1008 1456 2156 1512
rect 2352 1484 2772 1512
rect 2380 1456 2744 1484
rect 420 1428 700 1456
rect 476 1400 644 1428
rect 980 1400 2184 1456
rect 2464 1428 2688 1456
rect 952 1372 1512 1400
rect 1680 1372 2212 1400
rect 924 1344 1428 1372
rect 1764 1344 2240 1372
rect 924 1316 1372 1344
rect 1820 1316 2240 1344
rect 896 1288 1316 1316
rect 1876 1288 2268 1316
rect 868 1260 1288 1288
rect 1904 1260 2268 1288
rect 868 1232 1260 1260
rect 1932 1232 2296 1260
rect 840 1204 1232 1232
rect 812 1176 1232 1204
rect 1484 1176 1708 1204
rect 1960 1176 2324 1232
rect 812 1148 1204 1176
rect 1428 1148 1736 1176
rect 784 1092 1176 1148
rect 1400 1120 1764 1148
rect 1988 1120 2352 1176
rect 756 1064 1176 1092
rect 1372 1064 1792 1120
rect 2016 1064 2380 1120
rect 756 1036 1148 1064
rect 728 1008 1148 1036
rect 700 952 1148 1008
rect 672 896 1148 952
rect 1344 924 1820 1064
rect 2016 980 2408 1064
rect 2016 924 2436 980
rect 644 840 1176 896
rect 1372 868 1792 924
rect 2016 896 2464 924
rect 1988 868 2464 896
rect 1400 840 1764 868
rect 1988 840 2492 868
rect 616 812 1176 840
rect 1428 812 1736 840
rect 616 756 1204 812
rect 1484 784 1680 812
rect 1960 784 2492 840
rect 588 728 1232 756
rect 1932 728 2520 784
rect 588 700 1260 728
rect 1904 700 2548 728
rect 560 672 1288 700
rect 1876 672 2548 700
rect 560 644 1316 672
rect 1820 644 2548 672
rect 560 616 1372 644
rect 1792 616 2548 644
rect 532 588 1428 616
rect 1708 588 2576 616
rect 532 336 2576 588
rect 588 308 2520 336
<< end >>
