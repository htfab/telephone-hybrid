magic
tech sky130A
magscale 1 2
timestamp 1727597281
<< nwell >>
rect 0 954 48 2076
rect 2908 1952 2967 2010
rect 66 1078 124 1399
rect 2932 1078 2967 1952
rect 66 1020 148 1078
rect 2908 1020 2967 1078
rect 3008 954 3056 2076
<< pwell >>
rect 10 0 48 904
rect 2908 810 2926 868
rect 2908 36 2926 94
rect 3008 0 3056 904
<< mvpsubdiff >>
rect 46 810 148 868
rect 2908 810 3020 868
rect 46 760 104 810
rect 46 144 58 760
rect 92 144 104 760
rect 46 94 104 144
rect 2962 760 3020 810
rect 2962 144 2974 760
rect 3008 144 3020 760
rect 2962 94 3020 144
rect 46 36 148 94
rect 2908 36 3020 94
<< mvnsubdiff >>
rect 66 1952 148 2010
rect 2908 1952 2990 2010
rect 66 1902 124 1952
rect 66 1128 78 1902
rect 112 1128 124 1902
rect 66 1078 124 1128
rect 2932 1902 2990 1952
rect 2932 1128 2944 1902
rect 2978 1128 2990 1902
rect 2932 1078 2990 1128
rect 66 1020 148 1078
rect 2908 1020 2990 1078
<< mvpsubdiffcont >>
rect 58 144 92 760
rect 2974 144 3008 760
<< mvnsubdiffcont >>
rect 78 1128 112 1902
rect 2944 1128 2978 1902
<< locali >>
rect 78 1964 148 1998
rect 2908 1964 2978 1998
rect 78 1902 112 1964
rect 78 1066 112 1128
rect 2944 1902 2978 1964
rect 2944 1066 2978 1128
rect 78 1032 148 1066
rect 2908 1032 2978 1066
rect 58 822 148 856
rect 2908 822 3008 856
rect 58 760 92 822
rect 58 82 92 144
rect 2974 760 3008 822
rect 2974 82 3008 144
rect 58 48 148 82
rect 2908 48 3008 82
<< metal2 >>
rect 166 1866 2788 2004
rect 268 1193 406 1601
rect 2752 1193 2890 1601
rect 166 180 304 685
rect 452 557 570 675
rect 728 557 846 675
rect 1004 557 1122 675
rect 1280 557 1398 675
rect 1556 557 1674 675
rect 1832 557 1950 675
rect 2108 557 2226 675
rect 2384 557 2502 675
rect 2650 180 2788 685
rect 166 42 2788 180
<< via2 >>
rect 554 1203 672 1321
rect 830 1203 948 1321
rect 1106 1203 1224 1321
rect 1382 1203 1500 1321
rect 1658 1203 1776 1321
rect 1934 1203 2052 1321
rect 2210 1203 2328 1321
rect 2486 1203 2604 1321
<< metal3 >>
rect 544 1321 2614 1331
rect 544 1203 554 1321
rect 672 1203 830 1321
rect 948 1203 1106 1321
rect 1224 1203 1382 1321
rect 1500 1203 1658 1321
rect 1776 1203 1934 1321
rect 2052 1203 2210 1321
rect 2328 1203 2486 1321
rect 2604 1203 2614 1321
rect 544 1193 2614 1203
rect 622 1192 682 1193
rect 898 1192 958 1193
rect 1174 1192 1234 1193
rect 1450 1192 1510 1193
rect 1726 1192 1786 1193
rect 2002 1192 2062 1193
rect 2278 1192 2338 1193
rect 2554 1192 2614 1193
use passgate  x1
timestamp 1727597281
transform 1 0 324 0 1 0
box 0 0 476 2076
use passgate  x2
timestamp 1727597281
transform 1 0 600 0 1 0
box 0 0 476 2076
use passgate  x3
timestamp 1727597281
transform 1 0 876 0 1 0
box 0 0 476 2076
use passgate  x4
timestamp 1727597281
transform 1 0 1152 0 1 0
box 0 0 476 2076
use passgate  x5
timestamp 1727597281
transform 1 0 1428 0 1 0
box 0 0 476 2076
use passgate  x6
timestamp 1727597281
transform 1 0 1704 0 1 0
box 0 0 476 2076
use passgate  x7
timestamp 1727597281
transform 1 0 1980 0 1 0
box 0 0 476 2076
use passgate  x8
timestamp 1727597281
transform 1 0 2256 0 1 0
box 0 0 476 2076
use passgate  xdummy1
timestamp 1727597281
transform 1 0 48 0 1 0
box 0 0 476 2076
use passgate  xdummy2
timestamp 1727597281
transform 1 0 2532 0 1 0
box 0 0 476 2076
<< end >>
